
  --  Xilinx Single Port Byte-Write Read First RAM
  --  This code implements a parameterizable single-port byte-write read-first memory where when data
  --  is written to the memory, the output reflects the prior contents of the memory location.
  --  If a reset or enable is not necessary, it may be tied off or removed from the code.
  --  Modify the parameters for the desired RAM characteristics.

library ieee;
use ieee.std_logic_1164.all;

package ram_pkg is
    function clogb2 (depth: in natural) return integer;
end ram_pkg;

package body ram_pkg is

function clogb2( depth : natural) return integer is
variable temp    : integer := depth;
variable ret_val : integer := 0;
begin
    while temp > 1 loop
        ret_val := ret_val + 1;
        temp    := temp / 2;
   end loop;

   return ret_val;
end function;

end package body ram_pkg;

library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.ram_pkg.all;
USE std.textio.all;

entity RAM_Ins_48b is
--generic (
    --NB_COL    : integer;                       -- Specify number of columns (number of bytes)
    --COL_WIDTH : integer                       -- Specify column width (byte width, typically 8 or 9)
    --RAM_DEPTH : integer                        -- Specify RAM depth (number of entries)
 --   );

port (

        addra : in std_logic_vector(12 downto 0); 
        dina  : in std_logic_vector(47 downto 0);       -- RAM input data
        clka  : in std_logic;                           -- Clock
        wea   : in std_logic_vector(11 downto 0);        -- Byte-write enable
        ena   : in std_logic;                           -- RAM Enable, for additional power savings, disable port when not in use
        douta : out std_logic_vector(47 downto 0)       -- RAM output data
    );

end RAM_Ins_48b;

architecture rtl of RAM_Ins_48b is

constant C_NB_COL     : integer := 12;
constant C_COL_WIDTH  : integer := 4;
constant C_RAM_DEPTH  : integer := 8192; --512

signal douta_reg : std_logic_vector(C_NB_COL*C_COL_WIDTH-1 downto 0) := (others => '0');

--type ram_type is array (C_RAM_DEPTH-1 downto 0) of std_logic_vector (C_NB_COL*C_COL_WIDTH-1 downto 0);          -- 2D Array Declaration for RAM signal
type ram_type is array (0 to (C_RAM_DEPTH-1)) of std_logic_vector (C_NB_COL*C_COL_WIDTH-1 downto 0);  -- Modification necessaire pour remplir la mem � partir de l'adresse 0 C.JEGO 01/2025

signal ram_data : std_logic_vector(C_NB_COL*C_COL_WIDTH-1 downto 0) ;

--contenu de la m�moire instruction ; test consortium RISCV
signal ram_name : ram_type :=( X"00f300002537",
X"055f00050513",
X"0e5300450593",
X"0aac00b52023",
X"000300000093",
X"003f00000113",
X"003300000193",
X"005f00000213",
X"005300000293",
X"006f00000313",
X"006300000393",
X"006f00000413",
X"006300000493",
X"005f00000513",
X"005300000593",
X"003f00000613",
X"003300000693",
X"000f00000713",
X"000300000793",
X"007f00000813",
X"007300000893",
X"004f00000913",
X"004300000993",
X"002f00000a13",
X"002300000a93",
X"001f00000b13",
X"001300000b93",
X"001f00000c13",
X"001300000c93",
X"002f00000d13",
X"002300000d93",
X"004f00000e13",
X"004300000e93",
X"007f00000f13",
X"007300000f93",
X"20060a00006f",
X"0b063640006f",
X"79060810006f",
X"ae0627d0006f",
X"82067750006f",
X"f5067f90006f",
X"db962f40106f",
X"40966500106f",
X"d9961e10106f",
X"9e964dd0106f",
X"07a600c0206f",
X"10a63a00206f",
X"3ca63080206f",
X"a7a64cc0206f",
X"87a670c0206f",
X"fea614d0206f",
X"1ea63ad0206f",
X"49a66210206f",
X"0ea66bd0206f",
X"f73613c0306f",
X"6b363540306f",
X"52360550306f",
X"e2364250306f",
X"0cb60780406f",
X"4bb60940406f",
X"6bb63540406f",
X"49b60e10406f",
X"79b63910406f",
X"79b66410406f",
X"5b263440506f",
X"65260490506f",
X"5e2633d0506f",
X"ab161140606f",
X"40163f00606f",
X"89161b10606f",
X"3e166ad0606f",
X"00863100706f",
X"40865300706f",
X"000300000093",
X"00c100008067",
X"000300000093",
X"00cf00008713",
X"006300000393",
X"0a3300200193",
X"988726771c63",
X"090300100093",
X"09cf00108713",
X"0a6300200393",
X"033300300193",
X"98c726771263",
X"030300300093",
X"08cf00708713",
X"066300a00393",
X"0b3300400193",
X"c8e724771863",
X"000300000093",
X"c0cf80008713",
X"c06380000393",
X"023300500193",
X"f8d722771e63",
X"c00f800000b7",
X"00cf00008713",
X"c06f800003b7",
X"013300600193",
X"f8f722771463",
X"c00f800000b7",
X"c0cf80008713",
X"c06f800003b7",
X"c6a380038393",
X"083300700193",
X"a8e720771863",
X"000300000093",
X"f4cf7ff08713",
X"f4637ff00393",
X"0c3300800193",
X"d8d71e771e63",
X"c00f800000b7",
X"34c3fff08093",
X"00cf00008713",
X"c06f800003b7",
X"32a3fff38393",
X"053300900193",
X"d8971e771063",
X"c00f800000b7",
X"34c3fff08093",
X"f4cf7ff08713",
X"c06f800003b7",
X"fba37fe38393",
X"063300a00193",
X"88c71c771263",
X"c00f800000b7",
X"f4cf7ff08713",
X"c06f800003b7",
X"f2a37ff38393",
X"0f3300b00193",
X"b8a71a771663",
X"c00f800000b7",
X"34c3fff08093",
X"c0cf80008713",
X"f32f7ffff3b7",
X"f2a37ff38393",
X"073300c00193",
X"e8e718771863",
X"000300000093",
X"34cffff08713",
X"3463fff00393",
X"0e3300d00193",
X"a8d716771e63",
X"3403fff00093",
X"09cf00108713",
X"006300000393",
X"0d3300e00193",
X"a8f716771463",
X"3403fff00093",
X"34cffff08713",
X"3d63ffe00393",
X"043300f00193",
X"f8b714771a63",
X"c00f800000b7",
X"34c3fff08093",
X"09cf00108713",
X"c06f800003b7",
X"303301000193",
X"c8d712771e63",
X"0e0300d00093",
X"0fc300b08093",
X"3c6301800393",
X"393301100193",
X"c83712709463",
X"005f00000213",
X"0e0300d00093",
X"0fcf00b08713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"3c6301800393",
X"3a3301200193",
X"9e9710731063",
X"005f00000213",
X"0e0300d00093",
X"06cf00a08713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"386301700393",
X"333301300193",
X"1eb70c731a63",
X"005f00000213",
X"0e0300d00093",
X"05cf00908713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"316301600393",
X"3b3301400193",
X"2ec70a731263",
X"005f00000213",
X"0e0300d00093",
X"0fcf00b08713",
X"0c5f00120213",
X"0a5300200293",
X"07ebfe5218e3",
X"3c6301800393",
X"323301500193",
X"789708771063",
X"005f00000213",
X"0e0300d00093",
X"000f00000013",
X"06cf00a08713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"386301700393",
X"313301600193",
X"688704771c63",
X"005f00000213",
X"0e0300d00093",
X"000f00000013",
X"000f00000013",
X"05cf00908713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"316301600393",
X"383301700193",
X"58a702771663",
X"500302000093",
X"506302000393",
X"3c3301800193",
X"081700709e63",
X"590302100093",
X"6acf03208013",
X"006300000393",
X"353301900193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6e46cc1ff06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"5e46ca1ff06f",
X"000300000093",
X"003f00000113",
X"0ac500208733",
X"006300000393",
X"0a3300200193",
X"a8a74c771663",
X"090300100093",
X"093f00100113",
X"0ac500208733",
X"0a6300200393",
X"033300300193",
X"98b74a771a63",
X"030300300093",
X"083f00700113",
X"0ac500208733",
X"066300a00393",
X"0b3300400193",
X"c8d748771e63",
X"000300000093",
X"33f3ffff8137",
X"0ac500208733",
X"33afffff83b7",
X"023300500193",
X"c8c748771263",
X"c00f800000b7",
X"003f00000113",
X"0ac500208733",
X"c06f800003b7",
X"013300600193",
X"88a746771663",
X"c00f800000b7",
X"33f3ffff8137",
X"0ac500208733",
X"f3af7fff83b7",
X"083300700193",
X"d8b744771a63",
X"000300000093",
X"00f300008137",
X"373ffff10113",
X"0ac500208733",
X"00af000083b7",
X"32a3fff38393",
X"0c3300800193",
X"e8b742771a63",
X"c00f800000b7",
X"34c3fff08093",
X"003f00000113",
X"0ac500208733",
X"c06f800003b7",
X"32a3fff38393",
X"053300900193",
X"b8b740771a63",
X"c00f800000b7",
X"34c3fff08093",
X"00f300008137",
X"373ffff10113",
X"0ac500208733",
X"c0af800083b7",
X"3ba3ffe38393",
X"063300a00193",
X"78e73e771863",
X"c00f800000b7",
X"00f300008137",
X"373ffff10113",
X"0ac500208733",
X"c0af800083b7",
X"32a3fff38393",
X"0f3300b00193",
X"28e73c771863",
X"c00f800000b7",
X"34c3fff08093",
X"33f3ffff8137",
X"0ac500208733",
X"f3af7fff83b7",
X"32a3fff38393",
X"073300c00193",
X"18e73a771863",
X"000300000093",
X"343ffff00113",
X"0ac500208733",
X"3463fff00393",
X"0e3300d00193",
X"488738771c63",
X"3403fff00093",
X"093f00100113",
X"0ac500208733",
X"006300000393",
X"0d3300e00193",
X"489738771063",
X"3403fff00093",
X"343ffff00113",
X"0ac500208733",
X"3d63ffe00393",
X"043300f00193",
X"08f736771463",
X"090300100093",
X"c03380000137",
X"373ffff10113",
X"0ac500208733",
X"c06f800003b7",
X"303301000193",
X"58a734771663",
X"0e0300d00093",
X"0f3f00b00113",
X"0ac9002080b3",
X"3c6301800393",
X"393301100193",
X"687732709a63",
X"0d0300e00093",
X"0f3f00b00113",
X"0af500208133",
X"356301900393",
X"3a3301200193",
X"3bd730711e63",
X"0e0300d00093",
X"09c9001080b3",
X"366301a00393",
X"333301300193",
X"383730709463",
X"005f00000213",
X"0e0300d00093",
X"0f3f00b00113",
X"0ac500208733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"3c6301800393",
X"3b3301400193",
X"bed72c731e63",
X"005f00000213",
X"0d0300e00093",
X"0f3f00b00113",
X"0ac500208733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"356301900393",
X"323301500193",
X"8ea72a731663",
X"005f00000213",
X"040300f00093",
X"0f3f00b00113",
X"0ac500208733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"366301a00393",
X"313301600193",
X"9e8726731c63",
X"005f00000213",
X"0e0300d00093",
X"0f3f00b00113",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"3c6301800393",
X"383301700193",
X"c8e724771863",
X"005f00000213",
X"0d0300e00093",
X"0f3f00b00113",
X"000f00000013",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"356301900393",
X"3c3301800193",
X"f8c722771263",
X"005f00000213",
X"040300f00093",
X"0f3f00b00113",
X"000f00000013",
X"000f00000013",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"366301a00393",
X"353301900193",
X"d8b71e771a63",
X"005f00000213",
X"0e0300d00093",
X"000f00000013",
X"0f3f00b00113",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"3c6301800393",
X"363301a00193",
X"88f71c771463",
X"005f00000213",
X"0d0300e00093",
X"000f00000013",
X"0f3f00b00113",
X"000f00000013",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"356301900393",
X"3f3301b00193",
X"e88718771c63",
X"005f00000213",
X"040300f00093",
X"000f00000013",
X"000f00000013",
X"0f3f00b00113",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"366301a00393",
X"373301c00193",
X"a8f716771463",
X"005f00000213",
X"0f3f00b00113",
X"0e0300d00093",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"3c6301800393",
X"3e3301d00193",
X"f89714771063",
X"005f00000213",
X"0f3f00b00113",
X"0d0300e00093",
X"000f00000013",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"356301900393",
X"3d3301e00193",
X"98b710771a63",
X"005f00000213",
X"0f3f00b00113",
X"040300f00093",
X"000f00000013",
X"000f00000013",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"366301a00393",
X"343301f00193",
X"48c70e771263",
X"005f00000213",
X"0f3f00b00113",
X"000f00000013",
X"0e0300d00093",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"3c6301800393",
X"503302000193",
X"28870a771c63",
X"005f00000213",
X"0f3f00b00113",
X"000f00000013",
X"0d0300e00093",
X"000f00000013",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"356301900393",
X"593302100193",
X"78f708771463",
X"005f00000213",
X"0f3f00b00113",
X"000f00000013",
X"000f00000013",
X"040300f00093",
X"0ac500208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"366301a00393",
X"5a3302200193",
X"688704771c63",
X"040300f00093",
X"093500100133",
X"046300f00393",
X"533302300193",
X"6bc704711263",
X"500302000093",
X"00f500008133",
X"506302000393",
X"5b3302400193",
X"5be702711863",
X"0009000000b3",
X"006300000393",
X"523302500193",
X"585702709063",
X"300301000093",
X"3d3f01e00113",
X"0ac500208033",
X"006300000393",
X"513302600193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6c46fa4ff06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"3c46f84ff06f",
X"330fff0100b7",
X"40c3f0008093",
X"444ff0f0f713",
X"336fff0103b7",
X"46a3f0038393",
X"0a3300200193",
X"b8f71a771463",
X"749f0ff010b7",
X"30c3ff008093",
X"704f0f00f713",
X"70630f000393",
X"033300300193",
X"e8e718771863",
X"030f00ff00b7",
X"74c30ff08093",
X"844f70f0f713",
X"046300f00393",
X"0b3300400193",
X"a88716771c63",
X"474ff00ff0b7",
X"04c300f08093",
X"704f0f00f713",
X"006300000393",
X"023300500193",
X"a89716771063",
X"330fff0100b7",
X"40c3f0008093",
X"70430f00f093",
X"006300000393",
X"013300600193",
X"f83714709463",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"844f70f0f713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"806370000393",
X"083300700193",
X"9ed710731e63",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"704f0f00f713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"70630f000393",
X"0c3300800193",
X"4ea70e731663",
X"005f00000213",
X"474ff00ff0b7",
X"04c300f08093",
X"444ff0f0f713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"472ff00ff3b7",
X"02a300f38393",
X"053300900193",
X"2eb70a731a63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"844f70f0f713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"806370000393",
X"063300a00193",
X"78a708771663",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"704f0f00f713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"70630f000393",
X"0f3300b00193",
X"389706771063",
X"005f00000213",
X"474ff00ff0b7",
X"04c300f08093",
X"000f00000013",
X"000f00000013",
X"844f70f0f713",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"046300f00393",
X"073300c00193",
X"58e702771863",
X"70830f007093",
X"006300000393",
X"0e3300d00193",
X"585702709063",
X"030f00ff00b7",
X"74c30ff08093",
X"844f70f0f013",
X"006300000393",
X"0d3300e00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"cb46da8ff06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"9b46d88ff06f",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"70ff0f0013b7",
X"46a3f0038393",
X"0a3300200193",
X"c88748771c63",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0a450020f733",
X"046f00f003b7",
X"76a30f038393",
X"033300300193",
X"88b746771a63",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"076f000f03b7",
X"02a300f38393",
X"0b3300400193",
X"d8e744771863",
X"474ff00ff0b7",
X"04c300f08093",
X"4473f0f0f137",
X"733f0f010113",
X"0a450020f733",
X"402ff000f3b7",
X"023300500193",
X"e8e742771863",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a490020f0b3",
X"70ff0f0013b7",
X"46a3f0038393",
X"013300600193",
X"b86740709663",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0a750020f133",
X"046f00f003b7",
X"76a30f038393",
X"083300700193",
X"7bf73e711463",
X"330fff0100b7",
X"40c3f0008093",
X"09490010f0b3",
X"336fff0103b7",
X"46a3f0038393",
X"0c3300800193",
X"28673c709663",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"70ff0f0013b7",
X"46a3f0038393",
X"053300900193",
X"4eb738731a63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0a450020f733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"046f00f003b7",
X"76a30f038393",
X"063300a00193",
X"5e8734731c63",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"076f000f03b7",
X"02a300f38393",
X"0f3300b00193",
X"3e8730731c63",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"70ff0f0013b7",
X"46a3f0038393",
X"073300c00193",
X"e8c72e771263",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"046f00f003b7",
X"76a30f038393",
X"0e3300d00193",
X"88a72a771663",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"000f00000013",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"076f000f03b7",
X"02a300f38393",
X"0d3300e00193",
X"98e726771863",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"000f00000013",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"70ff0f0013b7",
X"46a3f0038393",
X"043300f00193",
X"f88722771c63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"046f00f003b7",
X"76a30f038393",
X"303301000193",
X"d8d71e771e63",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"000f00000013",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"076f000f03b7",
X"02a300f38393",
X"393301100193",
X"88971c771063",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"330fff0100b7",
X"40c3f0008093",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"70ff0f0013b7",
X"46a3f0038393",
X"3a3301200193",
X"e8a718771663",
X"005f00000213",
X"4473f0f0f137",
X"733f0f010113",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"046f00f003b7",
X"76a30f038393",
X"333301300193",
X"f8b714771a63",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"000f00000013",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"076f000f03b7",
X"02a300f38393",
X"3b3301400193",
X"988710771c63",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"330fff0100b7",
X"40c3f0008093",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"70ff0f0013b7",
X"46a3f0038393",
X"323301500193",
X"48970e771063",
X"005f00000213",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"046f00f003b7",
X"76a30f038393",
X"313301600193",
X"28c70a771263",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"000f00000013",
X"030f00ff00b7",
X"74c30ff08093",
X"0a450020f733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"076f000f03b7",
X"02a300f38393",
X"383301700193",
X"38f706771463",
X"330fff0100b7",
X"40c3f0008093",
X"09b500107133",
X"006300000393",
X"3c3301800193",
X"6be704711863",
X"030f00ff00b7",
X"74c30ff08093",
X"00750000f133",
X"006300000393",
X"353301900193",
X"5b8702711c63",
X"0089000070b3",
X"006300000393",
X"363301a00193",
X"583702709463",
X"aa9f111110b7",
X"a9c311108093",
X"ff9322222137",
X"f93f22210113",
X"0a450020f033",
X"006300000393",
X"3f3301b00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"dc468b4ff06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"8c46894ff06f",
X"000000000000",
X"00f900002517",
X"b25f71c50513",
X"0b5a004005ef",
X"ba5540b50533",
X"00cf000023b7",
X"b6a371038393",
X"0a3300200193",
X"5df702751463",
X"3389ffffe517",
X"b25f8fc50513",
X"0b5a004005ef",
X"ba5540b50533",
X"33bfffffe3b7",
X"b6a38f038393",
X"033300300193",
X"0df700751463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"a746830ff06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"f746810ff06f",
X"000000000000",
X"0a3300200193",
X"000300000093",
X"003f00000113",
X"0af700208663",
X"83e72a301863",
X"03a700301663",
X"0a8bfe208ee3",
X"83c72a301263",
X"033300300193",
X"090300100093",
X"093f00100113",
X"0af700208663",
X"d3e728301863",
X"03a700301663",
X"0a8bfe208ee3",
X"d3c728301263",
X"0b3300400193",
X"3403fff00093",
X"343ffff00113",
X"0af700208663",
X"93e726301863",
X"03a700301663",
X"0a8bfe208ee3",
X"93c726301263",
X"023300500193",
X"000300000093",
X"093f00100113",
X"0aa700208463",
X"03f700301463",
X"c3a724301663",
X"0a8bfe208ee3",
X"013300600193",
X"090300100093",
X"003f00000113",
X"0aa700208463",
X"03f700301463",
X"f3e722301863",
X"0a8bfe208ee3",
X"083300700193",
X"3403fff00093",
X"093f00100113",
X"0aa700208463",
X"03f700301463",
X"a3b720301a63",
X"0a8bfe208ee3",
X"0c3300800193",
X"090300100093",
X"343ffff00113",
X"0aa700208463",
X"03f700301463",
X"d3871e301c63",
X"0a8bfe208ee3",
X"053300900193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"dac71e208063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"063300a00193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"ba871a208e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0f3300b00193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"000f00000013",
X"eae718208a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"073300c00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"aab716208863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0e3300d00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"000f00000013",
X"faa714208463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0d3300e00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"343ffff00113",
X"cac712208063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"043300f00193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"9ac710208063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"303301000193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"1a870c208e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"393301100193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"000f00000013",
X"2ae70a208a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3a3301200193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"7ab708208863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"333301300193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"000f00000013",
X"3aa706208463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3b3301400193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"343ffff00113",
X"6ac704208063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"090300100093",
X"002700000a63",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"323301500193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"8ed6d31fe06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"ded6d11fe06f",
X"0a3300200193",
X"000300000093",
X"003f00000113",
X"0ad70020d663",
X"33e730301863",
X"03a700301663",
X"0aabfe20dee3",
X"33c730301263",
X"033300300193",
X"090300100093",
X"093f00100113",
X"0ad70020d663",
X"e3e72e301863",
X"03a700301663",
X"0aabfe20dee3",
X"e3c72e301263",
X"0b3300400193",
X"3403fff00093",
X"343ffff00113",
X"0ad70020d663",
X"b3e72c301863",
X"03a700301663",
X"0aabfe20dee3",
X"b3c72c301263",
X"023300500193",
X"090300100093",
X"003f00000113",
X"0ad70020d663",
X"83e72a301863",
X"03a700301663",
X"0aabfe20dee3",
X"83c72a301263",
X"013300600193",
X"090300100093",
X"343ffff00113",
X"0ad70020d663",
X"d3e728301863",
X"03a700301663",
X"0aabfe20dee3",
X"d3c728301263",
X"083300700193",
X"3403fff00093",
X"3d3fffe00113",
X"0ad70020d663",
X"93e726301863",
X"03a700301663",
X"0aabfe20dee3",
X"93c726301263",
X"0c3300800193",
X"000300000093",
X"093f00100113",
X"0a870020d463",
X"03f700301463",
X"c3a724301663",
X"0aabfe20dee3",
X"053300900193",
X"3403fff00093",
X"093f00100113",
X"0a870020d463",
X"03f700301463",
X"f3e722301863",
X"0aabfe20dee3",
X"063300a00193",
X"3d03ffe00093",
X"343ffff00113",
X"0a870020d463",
X"03f700301463",
X"a3b720301a63",
X"0aabfe20dee3",
X"0f3300b00193",
X"3d03ffe00093",
X"093f00100113",
X"0a870020d463",
X"03f700301463",
X"d3871e301c63",
X"0aabfe20dee3",
X"073300c00193",
X"005f00000213",
X"3403fff00093",
X"003f00000113",
X"dae71e20d063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"0e3300d00193",
X"005f00000213",
X"3403fff00093",
X"003f00000113",
X"000f00000013",
X"baa71a20de63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0d3300e00193",
X"005f00000213",
X"3403fff00093",
X"003f00000113",
X"000f00000013",
X"000f00000013",
X"eac71820da63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"043300f00193",
X"005f00000213",
X"3403fff00093",
X"000f00000013",
X"003f00000113",
X"aa971620d863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"303301000193",
X"005f00000213",
X"3403fff00093",
X"000f00000013",
X"003f00000113",
X"000f00000013",
X"fa871420d463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"393301100193",
X"005f00000213",
X"3403fff00093",
X"000f00000013",
X"000f00000013",
X"003f00000113",
X"cae71220d063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3a3301200193",
X"005f00000213",
X"3403fff00093",
X"003f00000113",
X"9ae71020d063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"333301300193",
X"005f00000213",
X"3403fff00093",
X"003f00000113",
X"000f00000013",
X"1aa70c20de63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"3b3301400193",
X"005f00000213",
X"3403fff00093",
X"003f00000113",
X"000f00000013",
X"000f00000013",
X"2ac70a20da63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"323301500193",
X"005f00000213",
X"3403fff00093",
X"000f00000013",
X"003f00000113",
X"7a970820d863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"313301600193",
X"005f00000213",
X"3403fff00093",
X"000f00000013",
X"003f00000113",
X"000f00000013",
X"3a870620d463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"383301700193",
X"005f00000213",
X"3403fff00093",
X"000f00000013",
X"000f00000013",
X"003f00000113",
X"6ae70420d063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"090300100093",
X"00c70000da63",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"3c3301800193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"75d69d5fe06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"45d69b5fe06f",
X"0a3300200193",
X"000300000093",
X"003f00000113",
X"0a770020f663",
X"53c734301263",
X"03a700301663",
X"0a0bfe20fee3",
X"638732301c63",
X"033300300193",
X"090300100093",
X"093f00100113",
X"0a770020f663",
X"63c732301263",
X"03a700301663",
X"0a0bfe20fee3",
X"338730301c63",
X"0b3300400193",
X"3403fff00093",
X"343ffff00113",
X"0a770020f663",
X"33c730301263",
X"03a700301663",
X"0a0bfe20fee3",
X"e3872e301c63",
X"023300500193",
X"090300100093",
X"003f00000113",
X"0a770020f663",
X"e3c72e301263",
X"03a700301663",
X"0a0bfe20fee3",
X"b3872c301c63",
X"013300600193",
X"3403fff00093",
X"3d3fffe00113",
X"0a770020f663",
X"b3c72c301263",
X"03a700301663",
X"0a0bfe20fee3",
X"83872a301c63",
X"083300700193",
X"3403fff00093",
X"003f00000113",
X"0a770020f663",
X"83c72a301263",
X"03a700301663",
X"0a0bfe20fee3",
X"d38728301c63",
X"0c3300800193",
X"000300000093",
X"093f00100113",
X"0a270020f463",
X"03f700301463",
X"d39728301063",
X"0a0bfe20fee3",
X"053300900193",
X"3d03ffe00093",
X"343ffff00113",
X"0a270020f463",
X"03f700301463",
X"93c726301263",
X"0a0bfe20fee3",
X"063300a00193",
X"000300000093",
X"343ffff00113",
X"0a270020f463",
X"03f700301463",
X"c3f724301463",
X"0a0bfe20fee3",
X"0f3300b00193",
X"c00f800000b7",
X"34c3fff08093",
X"c03380000137",
X"0a270020f463",
X"03f700301463",
X"f3f722301463",
X"0a0bfe20fee3",
X"073300c00193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"4033f0000137",
X"aa772020f663",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0e3300d00193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"4033f0000137",
X"000f00000013",
X"da171e20f263",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0d3300e00193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"4033f0000137",
X"000f00000013",
X"000f00000013",
X"ba571a20fc63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"043300f00193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"000f00000013",
X"4033f0000137",
X"ea371820f863",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"303301000193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"000f00000013",
X"4033f0000137",
X"000f00000013",
X"aa171620f263",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"393301100193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"000f00000013",
X"000f00000013",
X"4033f0000137",
X"ca571220fc63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"3a3301200193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"4033f0000137",
X"9a671020fa63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"333301300193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"4033f0000137",
X"000f00000013",
X"4a770e20f663",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3b3301400193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"4033f0000137",
X"000f00000013",
X"000f00000013",
X"1a470c20f063",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"323301500193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"000f00000013",
X"4033f0000137",
X"7a570820fc63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"313301600193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"000f00000013",
X"4033f0000137",
X"000f00000013",
X"3a770620f663",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"383301700193",
X"005f00000213",
X"400ff00000b7",
X"34c3fff08093",
X"000f00000013",
X"000f00000013",
X"4033f0000137",
X"6a470420f063",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"090300100093",
X"00670000fa63",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"3c3301800193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"bcd6e44fe06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"8cd6e24fe06f",
X"0a3300200193",
X"000300000093",
X"093f00100113",
X"0a470020c663",
X"83e72a301863",
X"03a700301663",
X"0a3bfe20cee3",
X"83c72a301263",
X"033300300193",
X"3403fff00093",
X"093f00100113",
X"0a470020c663",
X"d3e728301863",
X"03a700301663",
X"0a3bfe20cee3",
X"d3c728301263",
X"0b3300400193",
X"3d03ffe00093",
X"343ffff00113",
X"0a470020c663",
X"93e726301863",
X"03a700301663",
X"0a3bfe20cee3",
X"93c726301263",
X"023300500193",
X"090300100093",
X"003f00000113",
X"0a170020c463",
X"03f700301463",
X"c3a724301663",
X"0a3bfe20cee3",
X"013300600193",
X"090300100093",
X"343ffff00113",
X"0a170020c463",
X"03f700301463",
X"f3e722301863",
X"0a3bfe20cee3",
X"083300700193",
X"3403fff00093",
X"3d3fffe00113",
X"0a170020c463",
X"03f700301463",
X"a3b720301a63",
X"0a3bfe20cee3",
X"0c3300800193",
X"090300100093",
X"3d3fffe00113",
X"0a170020c463",
X"03f700301463",
X"d3871e301c63",
X"0a3bfe20cee3",
X"053300900193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"da771e20c063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"063300a00193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"ba371a20ce63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0f3300b00193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"000f00000013",
X"ea571820ca63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"073300c00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"aa071620c863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0e3300d00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"000f00000013",
X"fa171420c463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0d3300e00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"343ffff00113",
X"ca771220c063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"043300f00193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"9a771020c063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"303301000193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"1a370c20ce63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"393301100193",
X"005f00000213",
X"000300000093",
X"343ffff00113",
X"000f00000013",
X"000f00000013",
X"2a570a20ca63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3a3301200193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"7a070820c863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"333301300193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"343ffff00113",
X"000f00000013",
X"3a170620c463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3b3301400193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"343ffff00113",
X"6a770420c063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"090300100093",
X"099700104a63",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"323301500193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"9bd6b48fe06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"abd6b28fe06f",
X"0a3300200193",
X"000300000093",
X"093f00100113",
X"0ae70020e663",
X"e3c72e301263",
X"03a700301663",
X"0a9bfe20eee3",
X"b3872c301c63",
X"033300300193",
X"3d03ffe00093",
X"343ffff00113",
X"0ae70020e663",
X"b3c72c301263",
X"03a700301663",
X"0a9bfe20eee3",
X"83872a301c63",
X"0b3300400193",
X"000300000093",
X"343ffff00113",
X"0ae70020e663",
X"83c72a301263",
X"03a700301663",
X"0a9bfe20eee3",
X"d38728301c63",
X"023300500193",
X"090300100093",
X"003f00000113",
X"0ab70020e463",
X"03f700301463",
X"d39728301063",
X"0a9bfe20eee3",
X"013300600193",
X"3403fff00093",
X"3d3fffe00113",
X"0ab70020e463",
X"03f700301463",
X"93c726301263",
X"0a9bfe20eee3",
X"083300700193",
X"3403fff00093",
X"003f00000113",
X"0ab70020e463",
X"03f700301463",
X"c3f724301463",
X"0a9bfe20eee3",
X"0c3300800193",
X"c00f800000b7",
X"c03380000137",
X"373ffff10113",
X"0ab70020e463",
X"03f700301463",
X"f3f722301463",
X"0a9bfe20eee3",
X"053300900193",
X"005f00000213",
X"400ff00000b7",
X"4033f0000137",
X"373ffff10113",
X"aae72020e663",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"063300a00193",
X"005f00000213",
X"400ff00000b7",
X"4033f0000137",
X"373ffff10113",
X"000f00000013",
X"da871e20e263",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0f3300b00193",
X"005f00000213",
X"400ff00000b7",
X"4033f0000137",
X"373ffff10113",
X"000f00000013",
X"000f00000013",
X"bac71a20ec63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"073300c00193",
X"005f00000213",
X"400ff00000b7",
X"000f00000013",
X"4033f0000137",
X"373ffff10113",
X"eaa71820e863",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0e3300d00193",
X"005f00000213",
X"400ff00000b7",
X"000f00000013",
X"4033f0000137",
X"373ffff10113",
X"000f00000013",
X"aa871620e263",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0d3300e00193",
X"005f00000213",
X"400ff00000b7",
X"000f00000013",
X"000f00000013",
X"4033f0000137",
X"373ffff10113",
X"cac71220ec63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"043300f00193",
X"005f00000213",
X"400ff00000b7",
X"4033f0000137",
X"373ffff10113",
X"9af71020ea63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"303301000193",
X"005f00000213",
X"400ff00000b7",
X"4033f0000137",
X"373ffff10113",
X"000f00000013",
X"4ae70e20e663",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"393301100193",
X"005f00000213",
X"400ff00000b7",
X"4033f0000137",
X"373ffff10113",
X"000f00000013",
X"000f00000013",
X"1ad70c20e063",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"3a3301200193",
X"005f00000213",
X"400ff00000b7",
X"000f00000013",
X"4033f0000137",
X"373ffff10113",
X"7ac70820ec63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"333301300193",
X"005f00000213",
X"400ff00000b7",
X"000f00000013",
X"4033f0000137",
X"373ffff10113",
X"000f00000013",
X"3ae70620e663",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"3b3301400193",
X"005f00000213",
X"400ff00000b7",
X"000f00000013",
X"000f00000013",
X"4033f0000137",
X"373ffff10113",
X"6ad70420e063",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"090300100093",
X"093700106a63",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"323301500193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"fbd6818fe06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"32e6ff9fd06f",
X"0a3300200193",
X"000300000093",
X"093f00100113",
X"0a6700209663",
X"83b72a301a63",
X"03a700301663",
X"0a1bfe209ee3",
X"83f72a301463",
X"033300300193",
X"090300100093",
X"003f00000113",
X"0a6700209663",
X"d3b728301a63",
X"03a700301663",
X"0a1bfe209ee3",
X"d3f728301463",
X"0b3300400193",
X"3403fff00093",
X"093f00100113",
X"0a6700209663",
X"93b726301a63",
X"03a700301663",
X"0a1bfe209ee3",
X"93f726301463",
X"023300500193",
X"090300100093",
X"343ffff00113",
X"0a6700209663",
X"c3b724301a63",
X"03a700301663",
X"0a1bfe209ee3",
X"c3f724301463",
X"013300600193",
X"000300000093",
X"003f00000113",
X"0a3700209463",
X"03f700301463",
X"f3e722301863",
X"0a1bfe209ee3",
X"083300700193",
X"090300100093",
X"093f00100113",
X"0a3700209463",
X"03f700301463",
X"a3b720301a63",
X"0a1bfe209ee3",
X"0c3300800193",
X"3403fff00093",
X"343ffff00113",
X"0a3700209463",
X"03f700301463",
X"d3871e301c63",
X"0a1bfe209ee3",
X"053300900193",
X"005f00000213",
X"000300000093",
X"003f00000113",
X"da571e209063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"063300a00193",
X"005f00000213",
X"000300000093",
X"003f00000113",
X"000f00000013",
X"ba171a209e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0f3300b00193",
X"005f00000213",
X"000300000093",
X"003f00000113",
X"000f00000013",
X"000f00000013",
X"ea7718209a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"073300c00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"003f00000113",
X"aa2716209863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0e3300d00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"003f00000113",
X"000f00000013",
X"fa3714209463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0d3300e00193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"003f00000113",
X"ca5712209063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"043300f00193",
X"005f00000213",
X"000300000093",
X"003f00000113",
X"9a5710209063",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"303301000193",
X"005f00000213",
X"000300000093",
X"003f00000113",
X"000f00000013",
X"1a170c209e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"393301100193",
X"005f00000213",
X"000300000093",
X"003f00000113",
X"000f00000013",
X"000f00000013",
X"2a770a209a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3a3301200193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"003f00000113",
X"7a2708209863",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"333301300193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"003f00000113",
X"000f00000013",
X"3a3706209463",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3b3301400193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"003f00000113",
X"6a5704209063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"090300100093",
X"007700009a63",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"323301500193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"d2e6d19fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"02e6cf9fd06f",
X"0a3300200193",
X"000300000093",
X"30560100026f",
X"000f00000013",
X"000f00000013",
X"60060400006f",
X"003900000117",
X"383fff410113",
X"58b702411a63",
X"090300100093",
X"3b060140006f",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"09c300108093",
X"036300300393",
X"033300300193",
X"083700709463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"09e6c8dfd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"49e6c6dfd06f",
X"0a3300200193",
X"005300000293",
X"006900000317",
X"366f01030313",
X"065d000302e7",
X"40060e00006f",
X"006900000317",
X"316fffc30313",
X"14770c629a63",
X"033300300193",
X"005500000297",
X"359301028293",
X"059d000282e7",
X"10060c00006f",
X"006900000317",
X"316fffc30313",
X"24770a629a63",
X"0b3300400193",
X"005f00000213",
X"006900000317",
X"366f01030313",
X"063d000306e7",
X"73d708301e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"023300500193",
X"005f00000213",
X"006900000317",
X"3d6f01430313",
X"000f00000013",
X"063d000306e7",
X"33b706301a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"013300600193",
X"005f00000213",
X"006900000317",
X"3a6f01830313",
X"000f00000013",
X"000f00000013",
X"063d000306e7",
X"63f704301463",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"095300100293",
X"006900000317",
X"316f01c30313",
X"3101ffc30067",
X"0c9300128293",
X"0c9300128293",
X"0c9300128293",
X"0c9300128293",
X"0c9300128293",
X"0c9300128293",
X"0b6300400393",
X"083300700193",
X"0d3700729463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"a5e6b55fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"95e6b35fd06f",
X"000300000093",
X"00c600008703",
X"3463fff00393",
X"0a3300200193",
X"d8b71e771a63",
X"000300000093",
X"09c600108703",
X"006300000393",
X"033300300193",
X"d8971e771063",
X"000300000093",
X"0ac600208703",
X"3063ff000393",
X"0b3300400193",
X"88a71c771663",
X"000300000093",
X"03c600308703",
X"046300f00393",
X"023300500193",
X"b8871a771c63",
X"030300300093",
X"3ec6ffd08703",
X"3463fff00393",
X"013300600193",
X"b8c71a771263",
X"030300300093",
X"3dc6ffe08703",
X"006300000393",
X"083300700193",
X"e8e718771863",
X"030300300093",
X"34c6fff08703",
X"3063ff000393",
X"0c3300800193",
X"a8d716771e63",
X"030300300093",
X"00c600008703",
X"046300f00393",
X"053300900193",
X"a8f716771463",
X"000300000093",
X"00c3fe008093",
X"509a02008283",
X"3463fff00393",
X"063300a00193",
X"fd2714729863",
X"000300000093",
X"36c3ffa08093",
X"089a00708283",
X"006300000393",
X"0f3300b00193",
X"cd4712729c63",
X"073300c00193",
X"005f00000213",
X"090300100093",
X"09c600108703",
X"006f00070313",
X"3063ff000393",
X"9ed710731e63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0e3300d00193",
X"005f00000213",
X"0a0300200093",
X"09c600108703",
X"000f00000013",
X"006f00070313",
X"046300f00393",
X"4ee70e731863",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0d3300e00193",
X"005f00000213",
X"000300000093",
X"09c600108703",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"006300000393",
X"1e970c731063",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"043300f00193",
X"005f00000213",
X"090300100093",
X"09c600108703",
X"3063ff000393",
X"78d708771e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"303301000193",
X"005f00000213",
X"0a0300200093",
X"000f00000013",
X"09c600108703",
X"046300f00393",
X"38b706771a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"393301100193",
X"005f00000213",
X"000300000093",
X"000f00000013",
X"000f00000013",
X"09c600108703",
X"006300000393",
X"68f704771463",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"005300000293",
X"05f600028103",
X"0a3f00200113",
X"0a6300200393",
X"3a3301200193",
X"5bc702711263",
X"005300000293",
X"05f600028103",
X"000f00000013",
X"0a3f00200113",
X"0a6300200393",
X"333301300193",
X"0bf700711463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"62e6919fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"b2e68f9fd06f",
X"300301000093",
X"00760000c703",
X"74630ff00393",
X"0a3300200193",
X"d8b71e771a63",
X"300301000093",
X"09760010c703",
X"006300000393",
X"033300300193",
X"d8971e771063",
X"300301000093",
X"0a760020c703",
X"70630f000393",
X"0b3300400193",
X"88a71c771663",
X"300301000093",
X"03760030c703",
X"046300f00393",
X"023300500193",
X"b8871a771c63",
X"330301300093",
X"3e76ffd0c703",
X"74630ff00393",
X"013300600193",
X"b8c71a771263",
X"330301300093",
X"3d76ffe0c703",
X"006300000393",
X"083300700193",
X"e8e718771863",
X"330301300093",
X"3476fff0c703",
X"70630f000393",
X"0c3300800193",
X"a8d716771e63",
X"330301300093",
X"00760000c703",
X"046300f00393",
X"053300900193",
X"a8f716771463",
X"300301000093",
X"00c3fe008093",
X"502a0200c283",
X"74630ff00393",
X"063300a00193",
X"fd2714729863",
X"300301000093",
X"36c3ffa08093",
X"082a0070c283",
X"006300000393",
X"0f3300b00193",
X"cd4712729c63",
X"073300c00193",
X"005f00000213",
X"390301100093",
X"09760010c703",
X"006f00070313",
X"70630f000393",
X"9ed710731e63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0e3300d00193",
X"005f00000213",
X"3a0301200093",
X"09760010c703",
X"000f00000013",
X"006f00070313",
X"046300f00393",
X"4ee70e731863",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0d3300e00193",
X"005f00000213",
X"300301000093",
X"09760010c703",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"006300000393",
X"1e970c731063",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"043300f00193",
X"005f00000213",
X"390301100093",
X"09760010c703",
X"70630f000393",
X"78d708771e63",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"303301000193",
X"005f00000213",
X"3a0301200093",
X"000f00000013",
X"09760010c703",
X"046300f00393",
X"38b706771a63",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"393301100193",
X"005f00000213",
X"300301000093",
X"000f00000013",
X"000f00000013",
X"09760010c703",
X"006300000393",
X"68f704771463",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"305301000293",
X"05460002c103",
X"0a3f00200113",
X"0a6300200393",
X"3a3301200193",
X"5bc702711263",
X"305301000293",
X"05460002c103",
X"000f00000013",
X"0a3f00200113",
X"0a6300200393",
X"333301300193",
X"0bf700711463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"fbe6ed8fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"cbe6eb8fd06f",
X"500302000093",
X"005600009703",
X"74630ff00393",
X"0a3300200193",
X"a8b720771a63",
X"500302000093",
X"0a5600209703",
X"4063f0000393",
X"033300300193",
X"a89720771063",
X"500302000093",
X"0b5600409703",
X"00ff000013b7",
X"36a3ff038393",
X"0b3300400193",
X"d8f71e771463",
X"500302000093",
X"015600609703",
X"332ffffff3b7",
X"02a300f38393",
X"023300500193",
X"88e71c771863",
X"510302600093",
X"3656ffa09703",
X"74630ff00393",
X"013300600193",
X"b8d71a771e63",
X"510302600093",
X"3756ffc09703",
X"4063f0000393",
X"083300700193",
X"b8f71a771463",
X"510302600093",
X"3d56ffe09703",
X"00ff000013b7",
X"36a3ff038393",
X"0c3300800193",
X"e8e718771863",
X"510302600093",
X"005600009703",
X"332ffffff3b7",
X"02a300f38393",
X"053300900193",
X"a88716771c63",
X"500302000093",
X"00c3fe008093",
X"500a02009283",
X"74630ff00393",
X"063300a00193",
X"ad5716729063",
X"500302000093",
X"3fc3ffb08093",
X"080a00709283",
X"4063f0000393",
X"0f3300b00193",
X"fd3714729463",
X"073300c00193",
X"005f00000213",
X"5a0302200093",
X"0a5600209703",
X"006f00070313",
X"00ff000013b7",
X"36a3ff038393",
X"cef712731463",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0e3300d00193",
X"005f00000213",
X"5b0302400093",
X"0a5600209703",
X"000f00000013",
X"006f00070313",
X"332ffffff3b7",
X"02a300f38393",
X"4e870e731c63",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"0d3300e00193",
X"005f00000213",
X"500302000093",
X"0a5600209703",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"4063f0000393",
X"1ef70c731463",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"043300f00193",
X"005f00000213",
X"5a0302200093",
X"0a5600209703",
X"00ff000013b7",
X"36a3ff038393",
X"28970a771063",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"303301000193",
X"005f00000213",
X"5b0302400093",
X"000f00000013",
X"0a5600209703",
X"332ffffff3b7",
X"02a300f38393",
X"38b706771a63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"393301100193",
X"005f00000213",
X"500302000093",
X"000f00000013",
X"000f00000013",
X"0a5600209703",
X"4063f0000393",
X"68f704771463",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"505302000293",
X"056600029103",
X"0a3f00200113",
X"0a6300200393",
X"3a3301200193",
X"5bc702711263",
X"505302000293",
X"056600029103",
X"000f00000013",
X"0a3f00200113",
X"0a6300200393",
X"333301300193",
X"0bf700711463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"7be6c78fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"2be6c58fd06f",
X"600303000093",
X"00e60000d703",
X"74630ff00393",
X"0a3300200193",
X"f8f722771463",
X"600303000093",
X"0ae60020d703",
X"036f000103b7",
X"46a3f0038393",
X"033300300193",
X"a8e720771863",
X"600303000093",
X"0be60040d703",
X"00ff000013b7",
X"36a3ff038393",
X"0b3300400193",
X"d8871e771c63",
X"600303000093",
X"01e60060d703",
X"002f0000f3b7",
X"02a300f38393",
X"023300500193",
X"d8971e771063",
X"610303600093",
X"36e6ffa0d703",
X"74630ff00393",
X"013300600193",
X"88a71c771663",
X"610303600093",
X"37e6ffc0d703",
X"036f000103b7",
X"46a3f0038393",
X"083300700193",
X"b8b71a771a63",
X"610303600093",
X"3de6ffe0d703",
X"00ff000013b7",
X"36a3ff038393",
X"0c3300800193",
X"e8d718771e63",
X"610303600093",
X"00e60000d703",
X"002f0000f3b7",
X"02a300f38393",
X"053300900193",
X"e8c718771263",
X"600303000093",
X"00c3fe008093",
X"50ba0200d283",
X"74630ff00393",
X"063300a00193",
X"ad6716729663",
X"600303000093",
X"3fc3ffb08093",
X"08ba0070d283",
X"036f000103b7",
X"46a3f0038393",
X"0f3300b00193",
X"fd2714729863",
X"073300c00193",
X"005f00000213",
X"6a0303200093",
X"0ae60020d703",
X"006f00070313",
X"00ff000013b7",
X"36a3ff038393",
X"cee712731863",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0e3300d00193",
X"005f00000213",
X"6b0303400093",
X"0ae60020d703",
X"000f00000013",
X"006f00070313",
X"002f0000f3b7",
X"02a300f38393",
X"9e9710731063",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"0d3300e00193",
X"005f00000213",
X"600303000093",
X"0ae60020d703",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"036f000103b7",
X"46a3f0038393",
X"1ea70c731663",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"043300f00193",
X"005f00000213",
X"6a0303200093",
X"0ae60020d703",
X"00ff000013b7",
X"36a3ff038393",
X"28c70a771263",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"303301000193",
X"005f00000213",
X"6b0303400093",
X"000f00000013",
X"0ae60020d703",
X"002f0000f3b7",
X"02a300f38393",
X"388706771c63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"393301100193",
X"005f00000213",
X"600303000093",
X"000f00000013",
X"000f00000013",
X"0ae60020d703",
X"036f000103b7",
X"46a3f0038393",
X"68f704771463",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"605303000293",
X"05d60002d103",
X"0a3f00200113",
X"0a6300200393",
X"3a3301200193",
X"5bc702711263",
X"605303000293",
X"05d60002d103",
X"000f00000013",
X"0a3f00200113",
X"0a6300200393",
X"333301300193",
X"0bf700711463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6ce6a04fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"1ce69e4fd06f",
X"000f000000b7",
X"006300000393",
X"0a3300200193",
X"687704709a63",
X"334ffffff0b7",
X"b9e34010d093",
X"c06380000393",
X"033300300193",
X"685704709063",
X"f34f7ffff0b7",
X"8be34140d093",
X"f4637ff00393",
X"0b3300400193",
X"586702709663",
X"c00f800000b7",
X"8be34140d093",
X"c06380000393",
X"023300500193",
X"084700709c63",
X"c00380000037",
X"006300000393",
X"013300600193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6be6968fd06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"3be6948fd06f",
X"600304000093",
X"00660000a703",
X"036f00ff03b7",
X"72a30ff38393",
X"0a3300200193",
X"f8e722771863",
X"600304000093",
X"0b660040a703",
X"336fff0103b7",
X"46a3f0038393",
X"033300300193",
X"a88720771c63",
X"600304000093",
X"0c660080a703",
X"74ff0ff013b7",
X"36a3ff038393",
X"0b3300400193",
X"a89720771063",
X"600304000093",
X"076600c0a703",
X"472ff00ff3b7",
X"02a300f38393",
X"023300500193",
X"d8f71e771463",
X"670304c00093",
X"3b66ff40a703",
X"036f00ff03b7",
X"72a30ff38393",
X"013300600193",
X"88e71c771863",
X"670304c00093",
X"3c66ff80a703",
X"336fff0103b7",
X"46a3f0038393",
X"083300700193",
X"b8871a771c63",
X"670304c00093",
X"3766ffc0a703",
X"74ff0ff013b7",
X"36a3ff038393",
X"0c3300800193",
X"b8971a771063",
X"670304c00093",
X"00660000a703",
X"472ff00ff3b7",
X"02a300f38393",
X"053300900193",
X"e8f718771463",
X"600304000093",
X"00c3fe008093",
X"503a0200a283",
X"036f00ff03b7",
X"72a30ff38393",
X"063300a00193",
X"ad6716729663",
X"600304000093",
X"3ec3ffd08093",
X"083a0070a283",
X"336fff0103b7",
X"46a3f0038393",
X"0f3300b00193",
X"fd2714729863",
X"073300c00193",
X"005f00000213",
X"6b0304400093",
X"0b660040a703",
X"006f00070313",
X"74ff0ff013b7",
X"36a3ff038393",
X"cee712731863",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0e3300d00193",
X"005f00000213",
X"6c0304800093",
X"0b660040a703",
X"000f00000013",
X"006f00070313",
X"472ff00ff3b7",
X"02a300f38393",
X"9e9710731063",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"0d3300e00193",
X"005f00000213",
X"600304000093",
X"0b660040a703",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"336fff0103b7",
X"46a3f0038393",
X"1ea70c731663",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"043300f00193",
X"005f00000213",
X"6b0304400093",
X"0b660040a703",
X"74ff0ff013b7",
X"36a3ff038393",
X"28c70a771263",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"303301000193",
X"005f00000213",
X"6c0304800093",
X"000f00000013",
X"0b660040a703",
X"472ff00ff3b7",
X"02a300f38393",
X"388706771c63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"393301100193",
X"005f00000213",
X"600304000093",
X"000f00000013",
X"000f00000013",
X"0b660040a703",
X"336fff0103b7",
X"46a3f0038393",
X"68f704771463",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"605304000293",
X"05560002a103",
X"0a3f00200113",
X"0a6300200393",
X"3a3301200193",
X"5bc702711263",
X"605304000293",
X"05560002a103",
X"000f00000013",
X"0a3f00200113",
X"0a6300200393",
X"333301300193",
X"0bf700711463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"9276ee9fc06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"c276ec9fc06f",
X"330fff0100b7",
X"40c3f0008093",
X"44dff0f0e713",
X"4463f0f00393",
X"0a3300200193",
X"88f71c771463",
X"749f0ff010b7",
X"30c3ff008093",
X"70df0f00e713",
X"74ff0ff013b7",
X"36a3ff038393",
X"033300300193",
X"b8a71a771663",
X"030f00ff00b7",
X"74c30ff08093",
X"84df70f0e713",
X"036f00ff03b7",
X"f2a37ff38393",
X"0b3300400193",
X"e8e718771863",
X"474ff00ff0b7",
X"04c300f08093",
X"70df0f00e713",
X"472ff00ff3b7",
X"72a30ff38393",
X"023300500193",
X"a8b716771a63",
X"330fff0100b7",
X"40c3f0008093",
X"70d30f00e093",
X"336fff0103b7",
X"36a3ff038393",
X"013300600193",
X"f84714709c63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"70df0f00e713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"74ff0ff013b7",
X"36a3ff038393",
X"083300700193",
X"cef712731463",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"84df70f0e713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"036f00ff03b7",
X"f2a37ff38393",
X"0c3300800193",
X"4eb70e731a63",
X"005f00000213",
X"474ff00ff0b7",
X"04c300f08093",
X"70df0f00e713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"472ff00ff3b7",
X"72a30ff38393",
X"053300900193",
X"2ed70a731e63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"70df0f00e713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"74ff0ff013b7",
X"36a3ff038393",
X"063300a00193",
X"78e708771863",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"44dff0f0e713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"3463fff00393",
X"0f3300b00193",
X"38c706771263",
X"005f00000213",
X"474ff00ff0b7",
X"04c300f08093",
X"000f00000013",
X"000f00000013",
X"70df0f00e713",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"472ff00ff3b7",
X"72a30ff38393",
X"073300c00193",
X"58e702771863",
X"70130f006093",
X"70630f000393",
X"0e3300d00193",
X"585702709063",
X"030f00ff00b7",
X"74c30ff08093",
X"84df70f0e013",
X"006300000393",
X"0d3300e00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"5e76cd1fc06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6e76cb1fc06f",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"396fff1003b7",
X"42a3f0f38393",
X"0a3300200193",
X"98c74a771263",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0ad50020e733",
X"376ffff103b7",
X"36a3ff038393",
X"033300300193",
X"c89748771063",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"73ff0fff13b7",
X"32a3fff38393",
X"0b3300400193",
X"d8d744771e63",
X"474ff00ff0b7",
X"04c300f08093",
X"4473f0f0f137",
X"733f0f010113",
X"0ad50020e733",
X"432ff0fff3b7",
X"72a30ff38393",
X"023300500193",
X"e88742771c63",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad90020e0b3",
X"396fff1003b7",
X"42a3f0f38393",
X"013300600193",
X"b87740709a63",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ae50020e133",
X"396fff1003b7",
X"42a3f0f38393",
X"083300700193",
X"7be73e711863",
X"330fff0100b7",
X"40c3f0008093",
X"09d90010e0b3",
X"336fff0103b7",
X"46a3f0038393",
X"0c3300800193",
X"28773c709a63",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"396fff1003b7",
X"42a3f0f38393",
X"053300900193",
X"4ed738731e63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0ad50020e733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"376ffff103b7",
X"36a3ff038393",
X"063300a00193",
X"0e9736731063",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"73ff0fff13b7",
X"32a3fff38393",
X"0f3300b00193",
X"6e9732731063",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"396fff1003b7",
X"42a3f0f38393",
X"073300c00193",
X"e8a72e771663",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"376ffff103b7",
X"36a3ff038393",
X"0e3300d00193",
X"88b72a771a63",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"000f00000013",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"73ff0fff13b7",
X"32a3fff38393",
X"0d3300e00193",
X"988726771c63",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"000f00000013",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"396fff1003b7",
X"42a3f0f38393",
X"043300f00193",
X"c89724771063",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"376ffff103b7",
X"36a3ff038393",
X"303301000193",
X"a8c720771263",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"000f00000013",
X"77a30f0f1137",
X"473ff0f10113",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"73ff0fff13b7",
X"32a3fff38393",
X"393301100193",
X"88f71c771463",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"330fff0100b7",
X"40c3f0008093",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"396fff1003b7",
X"42a3f0f38393",
X"3a3301200193",
X"e8b718771a63",
X"005f00000213",
X"4473f0f0f137",
X"733f0f010113",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"376ffff103b7",
X"36a3ff038393",
X"333301300193",
X"f8d714771e63",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"000f00000013",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"73ff0fff13b7",
X"32a3fff38393",
X"3b3301400193",
X"c89712771063",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"330fff0100b7",
X"40c3f0008093",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"396fff1003b7",
X"42a3f0f38393",
X"323301500193",
X"48f70e771463",
X"005f00000213",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"376ffff103b7",
X"36a3ff038393",
X"313301600193",
X"28a70a771663",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"000f00000013",
X"030f00ff00b7",
X"74c30ff08093",
X"0ad50020e733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"73ff0fff13b7",
X"32a3fff38393",
X"383301700193",
X"38e706771863",
X"330fff0100b7",
X"40c3f0008093",
X"092500106133",
X"336fff0103b7",
X"46a3f0038393",
X"3c3301800193",
X"6bb704711a63",
X"030f00ff00b7",
X"74c30ff08093",
X"00e50000e133",
X"036f00ff03b7",
X"72a30ff38393",
X"353301900193",
X"5b8702711c63",
X"0019000060b3",
X"006300000393",
X"363301a00193",
X"583702709463",
X"aa9f111110b7",
X"a9c311108093",
X"ff9322222137",
X"f93f22210113",
X"0ad50020e033",
X"006300000393",
X"3f3301b00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6776fd0fc06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"5776fb0fc06f",
X"500305000093",
X"663ffaa00113",
X"0acc00208023",
X"00c600008703",
X"6663faa00393",
X"0a3300200193",
X"08d736771e63",
X"500305000093",
X"003f00000113",
X"0ac0002080a3",
X"09c600108703",
X"006300000393",
X"033300300193",
X"089736771063",
X"500305000093",
X"3373fffff137",
X"633ffa010113",
X"0afc00208123",
X"0a5600209703",
X"332ffffff3b7",
X"66a3fa038393",
X"0b3300400193",
X"68d732771e63",
X"500305000093",
X"063f00a00113",
X"0af0002081a3",
X"03c600308703",
X"066300a00393",
X"023300500193",
X"689732771063",
X"580305700093",
X"663ffaa00113",
X"0a80fe208ea3",
X"3ec6ffd08703",
X"6663faa00393",
X"013300600193",
X"38c730771263",
X"580305700093",
X"003f00000113",
X"0abcfe208f23",
X"3dc6ffe08703",
X"006300000393",
X"083300700193",
X"e8f72e771463",
X"580305700093",
X"603ffa000113",
X"0ab0fe208fa3",
X"34c6fff08703",
X"6063fa000393",
X"0c3300800193",
X"b8a72c771663",
X"580305700093",
X"063f00a00113",
X"0acc00208023",
X"00c600008703",
X"066300a00393",
X"053300900193",
X"88e72a771863",
X"5c0305800093",
X"c51312345137",
X"1f3f67810113",
X"009ffe008213",
X"5f0c02220023",
X"009a00008283",
X"0c6307800393",
X"063300a00193",
X"dd6728729663",
X"5c0305800093",
X"000300003137",
X"4f3f09810113",
X"36c3ffa08093",
X"0aa0002083a3",
X"555f05900213",
X"055a00020283",
X"0c63f9800393",
X"0f3300b00193",
X"9d0726729263",
X"073300c00193",
X"005f00000213",
X"6e03fdd00093",
X"503f05000113",
X"0a0c00110023",
X"030600010703",
X"6e63fdd00393",
X"c8c724771263",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0e3300d00193",
X"005f00000213",
X"5e03fcd00093",
X"503f05000113",
X"000f00000013",
X"0a00001100a3",
X"0a0600110703",
X"5e63fcd00393",
X"a8b720771a63",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"0d3300e00193",
X"005f00000213",
X"5703fcc00093",
X"503f05000113",
X"000f00000013",
X"000f00000013",
X"0a3c00110123",
X"090600210703",
X"5763fcc00393",
X"d8971e771063",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"043300f00193",
X"005f00000213",
X"5703fbc00093",
X"000f00000013",
X"503f05000113",
X"0a30001101a3",
X"000600310703",
X"5763fbc00393",
X"b8e71a771863",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"303301000193",
X"005f00000213",
X"5f03fbb00093",
X"000f00000013",
X"503f05000113",
X"000f00000013",
X"0a5c00110223",
X"080600410703",
X"5f63fbb00393",
X"a8d716771e63",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"393301100193",
X"005f00000213",
X"6f03fab00093",
X"000f00000013",
X"000f00000013",
X"503f05000113",
X"0a50001102a3",
X"010600510703",
X"6f63fab00393",
X"f8f714771463",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"3a3301200193",
X"005f00000213",
X"503f05000113",
X"630303300093",
X"0a0c00110023",
X"030600010703",
X"636303300393",
X"98d710771e63",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"333301300193",
X"005f00000213",
X"503f05000113",
X"530302300093",
X"000f00000013",
X"0a00001100a3",
X"0a0600110703",
X"536302300393",
X"48a70e771663",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"3b3301400193",
X"005f00000213",
X"503f05000113",
X"5a0302200093",
X"000f00000013",
X"000f00000013",
X"0a3c00110123",
X"090600210703",
X"5a6302200393",
X"28870a771c63",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"323301500193",
X"005f00000213",
X"503f05000113",
X"000f00000013",
X"3a0301200093",
X"0a30001101a3",
X"000600310703",
X"3a6301200393",
X"78f708771463",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"313301600193",
X"005f00000213",
X"503f05000113",
X"000f00000013",
X"390301100093",
X"000f00000013",
X"0a5c00110223",
X"080600410703",
X"396301100393",
X"68b704771a63",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"383301700193",
X"005f00000213",
X"503f05000113",
X"000f00000013",
X"000f00000013",
X"090300100093",
X"0a50001102a3",
X"010600510703",
X"096300100393",
X"589702771063",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"445f0ef00513",
X"505305000593",
X"03f000a581a3",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"7776c00fc06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"b776be0fc06f",
X"300306000093",
X"263f0aa00113",
X"0a5c00209023",
X"005600009703",
X"26630aa00393",
X"0a3300200193",
X"b89740771063",
X"300306000093",
X"33c3ffffb137",
X"633fa0010113",
X"0a6c00209123",
X"0a5600209703",
X"339fffffb3b7",
X"66a3a0038393",
X"033300300193",
X"28d73c771e63",
X"300306000093",
X"baa3beef1137",
X"433faa010113",
X"0a0c00209223",
X"0b660040a703",
X"baffbeef13b7",
X"46a3aa038393",
X"0b3300400193",
X"18873a771c63",
X"300306000093",
X"3353ffffa137",
X"053f00a10113",
X"0a3c00209323",
X"015600609703",
X"330fffffa3b7",
X"00a300a38393",
X"023300500193",
X"48b738771a63",
X"3d0306e00093",
X"263f0aa00113",
X"0a7cfe209d23",
X"3656ffa09703",
X"26630aa00393",
X"013300600193",
X"088736771c63",
X"3d0306e00093",
X"33c3ffffb137",
X"633fa0010113",
X"0a1cfe209e23",
X"3756ffc09703",
X"339fffffb3b7",
X"66a3a0038393",
X"083300700193",
X"58b734771a63",
X"3d0306e00093",
X"00a300001137",
X"433faa010113",
X"0a2cfe209f23",
X"3d56ffe09703",
X"00ff000013b7",
X"46a3aa038393",
X"0c3300800193",
X"68e732771863",
X"3d0306e00093",
X"3353ffffa137",
X"053f00a10113",
X"0a5c00209023",
X"005600009703",
X"330fffffa3b7",
X"00a300a38393",
X"053300900193",
X"38a730771663",
X"000307000093",
X"c51312345137",
X"1f3f67810113",
X"009ffe008213",
X"5f9c02221023",
X"000a00009283",
X"004f000053b7",
X"1aa367838393",
X"063300a00193",
X"ed072e729263",
X"000307000093",
X"000300003137",
X"4f3f09810113",
X"3fc3ffb08093",
X"0a30002093a3",
X"0a5f07200213",
X"05ca00021283",
X"005f000033b7",
X"4aa309838393",
X"0f3300b00193",
X"8d472a729c63",
X"073300c00193",
X"005f00000213",
X"33efffffd0b7",
X"5ec3cdd08093",
X"303f06000113",
X"0a9c00111023",
X"039600011703",
X"338fffffd3b7",
X"58a3cdd38393",
X"d8e728771863",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"0e3300d00193",
X"005f00000213",
X"337fffffc0b7",
X"6ec3ccd08093",
X"303f06000113",
X"000f00000013",
X"0aac00111123",
X"099600211703",
X"331fffffc3b7",
X"68a3ccd38393",
X"c88724771c63",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"0d3300e00193",
X"005f00000213",
X"337fffffc0b7",
X"e7c3bcc08093",
X"303f06000113",
X"000f00000013",
X"000f00000013",
X"0acc00111223",
X"089600411703",
X"331fffffc3b7",
X"e1a3bcc38393",
X"a8d720771e63",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"043300f00193",
X"005f00000213",
X"33ffffffb0b7",
X"e7c3bbc08093",
X"000f00000013",
X"303f06000113",
X"0afc00111323",
X"029600611703",
X"339fffffb3b7",
X"e1a3bbc38393",
X"d8c71e771263",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"303301000193",
X"005f00000213",
X"33ffffffb0b7",
X"7fc3abb08093",
X"000f00000013",
X"303f06000113",
X"000f00000013",
X"0afc00111423",
X"0f9600811703",
X"339fffffb3b7",
X"79a3abb38393",
X"b8f71a771463",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"393301100193",
X"005f00000213",
X"33dfffffe0b7",
X"4fc3aab08093",
X"000f00000013",
X"000f00000013",
X"303f06000113",
X"0acc00111523",
X"059600a11703",
X"33bfffffe3b7",
X"49a3aab38393",
X"a8a716771663",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"3a3301200193",
X"005f00000213",
X"303f06000113",
X"00af000020b7",
X"c3c323308093",
X"0a9c00111023",
X"039600011703",
X"00cf000023b7",
X"c5a323338393",
X"c88712771c63",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"333301300193",
X"005f00000213",
X"303f06000113",
X"009f000010b7",
X"f3c322308093",
X"000f00000013",
X"0aac00111123",
X"099600211703",
X"00ff000013b7",
X"f5a322338393",
X"989710771063",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"3b3301400193",
X"005f00000213",
X"303f06000113",
X"009f000010b7",
X"cac312208093",
X"000f00000013",
X"000f00000013",
X"0acc00111223",
X"089600411703",
X"00ff000013b7",
X"cca312238393",
X"18c70c771263",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"323301500193",
X"005f00000213",
X"303f06000113",
X"000f00000013",
X"aa0311200093",
X"0afc00111323",
X"029600611703",
X"aa6311200393",
X"78b708771a63",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"313301600193",
X"005f00000213",
X"303f06000113",
X"000f00000013",
X"390301100093",
X"000f00000013",
X"0afc00111423",
X"0f9600811703",
X"396301100393",
X"389706771063",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"383301700193",
X"005f00000213",
X"303f06000113",
X"000f00000013",
X"000f00000013",
X"003f000030b7",
X"09c300108093",
X"0acc00111523",
X"059600a11703",
X"005f000033b7",
X"0fa300138393",
X"58c702771263",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"00230000c537",
X"915feef50513",
X"305306000593",
X"033c00a59323",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"69f6fadfb06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"39f6f8dfb06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"4ef6f71fb06f",
X"090300100093",
X"005f00009713",
X"096300100393",
X"0a3300200193",
X"98b726771a63",
X"090300100093",
X"095f00109713",
X"0a6300200393",
X"033300300193",
X"989726771063",
X"090300100093",
X"085f00709713",
X"706308000393",
X"0b3300400193",
X"c8a724771663",
X"090300100093",
X"0d5f00e09713",
X"00df000043b7",
X"023300500193",
X"f88722771c63",
X"090300100093",
X"345f01f09713",
X"c06f800003b7",
X"013300600193",
X"f8c722771263",
X"3403fff00093",
X"005f00009713",
X"3463fff00393",
X"083300700193",
X"a8e720771863",
X"3403fff00093",
X"095f00109713",
X"3d63ffe00393",
X"0c3300800193",
X"d8d71e771e63",
X"3403fff00093",
X"085f00709713",
X"3063f8000393",
X"053300900193",
X"d8f71e771463",
X"3403fff00093",
X"0d5f00e09713",
X"331fffffc3b7",
X"063300a00193",
X"88b71c771a63",
X"3403fff00093",
X"345f01f09713",
X"c06f800003b7",
X"0f3300b00193",
X"88971c771063",
X"99af212120b7",
X"c9c312108093",
X"005f00009713",
X"99cf212123b7",
X"cfa312138393",
X"073300c00193",
X"b8c71a771263",
X"99af212120b7",
X"c9c312108093",
X"095f00109713",
X"eedf424243b7",
X"cca324238393",
X"0e3300d00193",
X"e8f718771463",
X"99af212120b7",
X"c9c312108093",
X"085f00709713",
X"553f909093b7",
X"76a308038393",
X"0d3300e00193",
X"a8a716771663",
X"99af212120b7",
X"c9c312108093",
X"0d5f00e09713",
X"ccdf484843b7",
X"043300f00193",
X"f8b714771a63",
X"99af212120b7",
X"c9c312108093",
X"345f01f09713",
X"c06f800003b7",
X"303301000193",
X"c8d712771e63",
X"090300100093",
X"085300709093",
X"706308000393",
X"393301100193",
X"c83712709463",
X"005f00000213",
X"090300100093",
X"085f00709713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"706308000393",
X"3a3301200193",
X"9e9710731063",
X"005f00000213",
X"090300100093",
X"0d5f00e09713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"00df000043b7",
X"333301300193",
X"1eb70c731a63",
X"005f00000213",
X"090300100093",
X"345f01f09713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"c06f800003b7",
X"3b3301400193",
X"2ec70a731263",
X"005f00000213",
X"090300100093",
X"085f00709713",
X"0c5f00120213",
X"0a5300200293",
X"07ebfe5218e3",
X"706308000393",
X"323301500193",
X"789708771063",
X"005f00000213",
X"090300100093",
X"000f00000013",
X"0d5f00e09713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"00df000043b7",
X"313301600193",
X"688704771c63",
X"005f00000213",
X"090300100093",
X"000f00000013",
X"000f00000013",
X"345f01f09713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"c06f800003b7",
X"383301700193",
X"58a702771663",
X"349301f01093",
X"006300000393",
X"3c3301800193",
X"081700709e63",
X"590302100093",
X"3b5f01409013",
X"006300000393",
X"353301900193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"5ef6cd1fb06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6ef6cb1fb06f",
X"090300100093",
X"003f00000113",
X"0a5500209733",
X"096300100393",
X"0a3300200193",
X"78d752771e63",
X"090300100093",
X"093f00100113",
X"0a5500209733",
X"0a6300200393",
X"033300300193",
X"78c752771263",
X"090300100093",
X"083f00700113",
X"0a5500209733",
X"706308000393",
X"0b3300400193",
X"28a750771663",
X"090300100093",
X"0d3f00e00113",
X"0a5500209733",
X"00df000043b7",
X"023300500193",
X"f8b74e771a63",
X"090300100093",
X"343f01f00113",
X"0a5500209733",
X"c06f800003b7",
X"013300600193",
X"a8d74c771e63",
X"3403fff00093",
X"003f00000113",
X"0a5500209733",
X"3463fff00393",
X"083300700193",
X"a8c74c771263",
X"3403fff00093",
X"093f00100113",
X"0a5500209733",
X"3d63ffe00393",
X"0c3300800193",
X"98a74a771663",
X"3403fff00093",
X"083f00700113",
X"0a5500209733",
X"3063f8000393",
X"053300900193",
X"c8b748771a63",
X"3403fff00093",
X"0d3f00e00113",
X"0a5500209733",
X"331fffffc3b7",
X"063300a00193",
X"88d746771e63",
X"3403fff00093",
X"343f01f00113",
X"0a5500209733",
X"c06f800003b7",
X"0f3300b00193",
X"88c746771263",
X"99af212120b7",
X"c9c312108093",
X"003f00000113",
X"0a5500209733",
X"99cf212123b7",
X"cfa312138393",
X"073300c00193",
X"d8c744771263",
X"99af212120b7",
X"c9c312108093",
X"093f00100113",
X"0a5500209733",
X"eedf424243b7",
X"cca324238393",
X"0e3300d00193",
X"e8c742771263",
X"99af212120b7",
X"c9c312108093",
X"083f00700113",
X"0a5500209733",
X"553f909093b7",
X"76a308038393",
X"0d3300e00193",
X"b8c740771263",
X"99af212120b7",
X"c9c312108093",
X"0d3f00e00113",
X"0a5500209733",
X"ccdf484843b7",
X"043300f00193",
X"78f73e771463",
X"99af212120b7",
X"c9c312108093",
X"343f01f00113",
X"0a5500209733",
X"c06f800003b7",
X"303301000193",
X"28a73c771663",
X"99af212120b7",
X"c9c312108093",
X"503ffc000113",
X"0a5500209733",
X"99cf212123b7",
X"cfa312138393",
X"393301100193",
X"18a73a771663",
X"99af212120b7",
X"c9c312108093",
X"593ffc100113",
X"0a5500209733",
X"eedf424243b7",
X"cca324238393",
X"3a3301200193",
X"48a738771663",
X"99af212120b7",
X"c9c312108093",
X"583ffc700113",
X"0a5500209733",
X"553f909093b7",
X"76a308038393",
X"333301300193",
X"08a736771663",
X"99af212120b7",
X"c9c312108093",
X"5d3ffce00113",
X"0a5500209733",
X"ccdf484843b7",
X"3b3301400193",
X"58e734771863",
X"090300100093",
X"083f00700113",
X"0a59002090b3",
X"706308000393",
X"313301600193",
X"684732709c63",
X"090300100093",
X"0d3f00e00113",
X"0a6500209133",
X"00df000043b7",
X"383301700193",
X"6b9732711063",
X"030300300093",
X"0959001090b3",
X"3c6301800393",
X"3c3301800193",
X"386730709663",
X"005f00000213",
X"090300100093",
X"083f00700113",
X"0a5500209733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"706308000393",
X"353301900193",
X"ee972e731063",
X"005f00000213",
X"090300100093",
X"0d3f00e00113",
X"0a5500209733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"00df000043b7",
X"363301a00193",
X"8ee72a731863",
X"005f00000213",
X"090300100093",
X"343f01f00113",
X"0a5500209733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"c06f800003b7",
X"3f3301b00193",
X"9ed726731e63",
X"005f00000213",
X"090300100093",
X"083f00700113",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"706308000393",
X"373301c00193",
X"c8b724771a63",
X"005f00000213",
X"090300100093",
X"0d3f00e00113",
X"000f00000013",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"00df000043b7",
X"3e3301d00193",
X"f8f722771463",
X"005f00000213",
X"090300100093",
X"343f01f00113",
X"000f00000013",
X"000f00000013",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"c06f800003b7",
X"3d3301e00193",
X"d8871e771c63",
X"005f00000213",
X"090300100093",
X"000f00000013",
X"083f00700113",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"706308000393",
X"343301f00193",
X"88a71c771663",
X"005f00000213",
X"090300100093",
X"000f00000013",
X"0d3f00e00113",
X"000f00000013",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"00df000043b7",
X"503302000193",
X"e8d718771e63",
X"005f00000213",
X"090300100093",
X"000f00000013",
X"000f00000013",
X"343f01f00113",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"c06f800003b7",
X"593302100193",
X"a8a716771663",
X"005f00000213",
X"083f00700113",
X"090300100093",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"706308000393",
X"5a3302200193",
X"f8c714771263",
X"005f00000213",
X"0d3f00e00113",
X"090300100093",
X"000f00000013",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"00df000043b7",
X"533302300193",
X"988710771c63",
X"005f00000213",
X"343f01f00113",
X"090300100093",
X"000f00000013",
X"000f00000013",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"c06f800003b7",
X"5b3302400193",
X"48f70e771463",
X"005f00000213",
X"083f00700113",
X"000f00000013",
X"090300100093",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"706308000393",
X"523302500193",
X"28d70a771e63",
X"005f00000213",
X"0d3f00e00113",
X"000f00000013",
X"090300100093",
X"000f00000013",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"00df000043b7",
X"513302600193",
X"78a708771663",
X"005f00000213",
X"343f01f00113",
X"000f00000013",
X"000f00000013",
X"090300100093",
X"0a5500209733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"c06f800003b7",
X"583302700193",
X"68d704771e63",
X"040300f00093",
X"09a500101133",
X"006300000393",
X"5c3302800193",
X"6bf704711463",
X"500302000093",
X"006500009133",
X"506302000393",
X"553302900193",
X"5bb702711a63",
X"0099000010b3",
X"006300000393",
X"563302a00193",
X"580702709263",
X"b00340000093",
X"00a300001137",
X"c33f80010113",
X"0a5500209033",
X"006300000393",
X"5f3302b00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"2cf6f44fb06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"1cf6f24fb06f",
X"000300000093",
X"006f0000a713",
X"006300000393",
X"0a3300200193",
X"98c726771263",
X"090300100093",
X"096f0010a713",
X"006300000393",
X"033300300193",
X"c8e724771863",
X"030300300093",
X"086f0070a713",
X"096300100393",
X"0b3300400193",
X"f8d722771e63",
X"080300700093",
X"036f0030a713",
X"006300000393",
X"023300500193",
X"f8f722771463",
X"000300000093",
X"c06f8000a713",
X"006300000393",
X"013300600193",
X"a8b720771a63",
X"c00f800000b7",
X"006f0000a713",
X"096300100393",
X"083300700193",
X"a89720771063",
X"c00f800000b7",
X"c06f8000a713",
X"096300100393",
X"0c3300800193",
X"d8a71e771663",
X"000300000093",
X"f46f7ff0a713",
X"096300100393",
X"053300900193",
X"88871c771c63",
X"c00f800000b7",
X"34c3fff08093",
X"006f0000a713",
X"006300000393",
X"063300a00193",
X"88971c771063",
X"c00f800000b7",
X"34c3fff08093",
X"f46f7ff0a713",
X"006300000393",
X"0f3300b00193",
X"b8f71a771463",
X"c00f800000b7",
X"f46f7ff0a713",
X"096300100393",
X"073300c00193",
X"e8b718771a63",
X"c00f800000b7",
X"34c3fff08093",
X"c06f8000a713",
X"006300000393",
X"0e3300d00193",
X"a8d716771e63",
X"000300000093",
X"346ffff0a713",
X"006300000393",
X"0d3300e00193",
X"a8f716771463",
X"3403fff00093",
X"096f0010a713",
X"096300100393",
X"043300f00193",
X"f8b714771a63",
X"3403fff00093",
X"346ffff0a713",
X"006300000393",
X"303301000193",
X"f89714771063",
X"0f0300b00093",
X"0e6300d0a093",
X"096300100393",
X"393301100193",
X"c86712709663",
X"005f00000213",
X"040300f00093",
X"066f00a0a713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"3a3301200193",
X"9ec710731263",
X"005f00000213",
X"060300a00093",
X"306f0100a713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"333301300193",
X"1e870c731c63",
X"005f00000213",
X"300301000093",
X"056f0090a713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"3b3301400193",
X"2ef70a731463",
X"005f00000213",
X"0f0300b00093",
X"046f00f0a713",
X"0c5f00120213",
X"0a5300200293",
X"07ebfe5218e3",
X"096300100393",
X"323301500193",
X"78c708771263",
X"005f00000213",
X"390301100093",
X"000f00000013",
X"0c6f0080a713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"313301600193",
X"68d704771e63",
X"005f00000213",
X"070300c00093",
X"000f00000013",
X"000f00000013",
X"0d6f00e0a713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"383301700193",
X"58e702771863",
X"34a3fff02093",
X"006300000393",
X"3c3301800193",
X"585702709063",
X"030f00ff00b7",
X"74c30ff08093",
X"346ffff0a013",
X"006300000393",
X"353301900193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"3cf6c94fb06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"7cf6c74fb06f",
X"000300000093",
X"00ff0000b713",
X"006300000393",
X"0a3300200193",
X"98c726771263",
X"090300100093",
X"09ff0010b713",
X"006300000393",
X"033300300193",
X"c8e724771863",
X"030300300093",
X"08ff0070b713",
X"096300100393",
X"0b3300400193",
X"f8d722771e63",
X"080300700093",
X"03ff0030b713",
X"006300000393",
X"023300500193",
X"f8f722771463",
X"000300000093",
X"c0ff8000b713",
X"096300100393",
X"013300600193",
X"a8b720771a63",
X"c00f800000b7",
X"00ff0000b713",
X"006300000393",
X"083300700193",
X"a89720771063",
X"c00f800000b7",
X"c0ff8000b713",
X"096300100393",
X"0c3300800193",
X"d8a71e771663",
X"000300000093",
X"f4ff7ff0b713",
X"096300100393",
X"053300900193",
X"88871c771c63",
X"c00f800000b7",
X"34c3fff08093",
X"00ff0000b713",
X"006300000393",
X"063300a00193",
X"88971c771063",
X"c00f800000b7",
X"34c3fff08093",
X"f4ff7ff0b713",
X"006300000393",
X"0f3300b00193",
X"b8f71a771463",
X"c00f800000b7",
X"f4ff7ff0b713",
X"006300000393",
X"073300c00193",
X"e8b718771a63",
X"c00f800000b7",
X"34c3fff08093",
X"c0ff8000b713",
X"096300100393",
X"0e3300d00193",
X"a8d716771e63",
X"000300000093",
X"34fffff0b713",
X"096300100393",
X"0d3300e00193",
X"a8f716771463",
X"3403fff00093",
X"09ff0010b713",
X"006300000393",
X"043300f00193",
X"f8b714771a63",
X"3403fff00093",
X"34fffff0b713",
X"006300000393",
X"303301000193",
X"f89714771063",
X"0f0300b00093",
X"0ef300d0b093",
X"096300100393",
X"393301100193",
X"c86712709663",
X"005f00000213",
X"040300f00093",
X"06ff00a0b713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"3a3301200193",
X"9ec710731263",
X"005f00000213",
X"060300a00093",
X"30ff0100b713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"333301300193",
X"1e870c731c63",
X"005f00000213",
X"300301000093",
X"05ff0090b713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"3b3301400193",
X"2ef70a731463",
X"005f00000213",
X"0f0300b00093",
X"04ff00f0b713",
X"0c5f00120213",
X"0a5300200293",
X"07ebfe5218e3",
X"096300100393",
X"323301500193",
X"78c708771263",
X"005f00000213",
X"390301100093",
X"000f00000013",
X"0cff0080b713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"313301600193",
X"68d704771e63",
X"005f00000213",
X"070300c00093",
X"000f00000013",
X"000f00000013",
X"0dff00e0b713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"383301700193",
X"58e702771863",
X"3433fff03093",
X"096300100393",
X"3c3301800193",
X"585702709063",
X"030f00ff00b7",
X"74c30ff08093",
X"34fffff0b013",
X"006300000393",
X"353301900193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"1cf69e4fb06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"4cf69c4fb06f",
X"000300000093",
X"003f00000113",
X"0a650020a733",
X"006300000393",
X"0a3300200193",
X"98b74a771a63",
X"090300100093",
X"093f00100113",
X"0a650020a733",
X"006300000393",
X"033300300193",
X"c8d748771e63",
X"030300300093",
X"083f00700113",
X"0a650020a733",
X"096300100393",
X"0b3300400193",
X"c8c748771263",
X"080300700093",
X"033f00300113",
X"0a650020a733",
X"006300000393",
X"023300500193",
X"88a746771663",
X"000300000093",
X"33f3ffff8137",
X"0a650020a733",
X"006300000393",
X"013300600193",
X"d8b744771a63",
X"c00f800000b7",
X"003f00000113",
X"0a650020a733",
X"096300100393",
X"083300700193",
X"e8d742771e63",
X"c00f800000b7",
X"33f3ffff8137",
X"0a650020a733",
X"096300100393",
X"0c3300800193",
X"e8c742771263",
X"000300000093",
X"00f300008137",
X"373ffff10113",
X"0a650020a733",
X"096300100393",
X"053300900193",
X"b8f740771463",
X"c00f800000b7",
X"34c3fff08093",
X"003f00000113",
X"0a650020a733",
X"006300000393",
X"063300a00193",
X"78a73e771663",
X"c00f800000b7",
X"34c3fff08093",
X"00f300008137",
X"373ffff10113",
X"0a650020a733",
X"006300000393",
X"0f3300b00193",
X"28a73c771663",
X"c00f800000b7",
X"00f300008137",
X"373ffff10113",
X"0a650020a733",
X"096300100393",
X"073300c00193",
X"18e73a771863",
X"c00f800000b7",
X"34c3fff08093",
X"33f3ffff8137",
X"0a650020a733",
X"006300000393",
X"0e3300d00193",
X"48b738771a63",
X"000300000093",
X"343ffff00113",
X"0a650020a733",
X"006300000393",
X"0d3300e00193",
X"08d736771e63",
X"3403fff00093",
X"093f00100113",
X"0a650020a733",
X"096300100393",
X"043300f00193",
X"08c736771263",
X"3403fff00093",
X"343ffff00113",
X"0a650020a733",
X"006300000393",
X"303301000193",
X"58a734771663",
X"0d0300e00093",
X"0e3f00d00113",
X"0a690020a0b3",
X"006300000393",
X"393301100193",
X"687732709a63",
X"0f0300b00093",
X"0e3f00d00113",
X"0a550020a133",
X"096300100393",
X"3a3301200193",
X"3bd730711e63",
X"0e0300d00093",
X"09690010a0b3",
X"006300000393",
X"333301300193",
X"383730709463",
X"005f00000213",
X"0f0300b00093",
X"0e3f00d00113",
X"0a650020a733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"3b3301400193",
X"bed72c731e63",
X"005f00000213",
X"0d0300e00093",
X"0e3f00d00113",
X"0a650020a733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"323301500193",
X"8ea72a731663",
X"005f00000213",
X"070300c00093",
X"0e3f00d00113",
X"0a650020a733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"096300100393",
X"313301600193",
X"9e8726731c63",
X"005f00000213",
X"0d0300e00093",
X"0e3f00d00113",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"383301700193",
X"c8e724771863",
X"005f00000213",
X"0f0300b00093",
X"0e3f00d00113",
X"000f00000013",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"3c3301800193",
X"f8c722771263",
X"005f00000213",
X"040300f00093",
X"0e3f00d00113",
X"000f00000013",
X"000f00000013",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"353301900193",
X"d8b71e771a63",
X"005f00000213",
X"060300a00093",
X"000f00000013",
X"0e3f00d00113",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"363301a00193",
X"88f71c771463",
X"005f00000213",
X"300301000093",
X"000f00000013",
X"0e3f00d00113",
X"000f00000013",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"3f3301b00193",
X"e88718771c63",
X"005f00000213",
X"050300900093",
X"000f00000013",
X"000f00000013",
X"0e3f00d00113",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"373301c00193",
X"a8f716771463",
X"005f00000213",
X"0e3f00d00113",
X"390301100093",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"3e3301d00193",
X"f89714771063",
X"005f00000213",
X"0e3f00d00113",
X"0c0300800093",
X"000f00000013",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"3d3301e00193",
X"98b710771a63",
X"005f00000213",
X"0e3f00d00113",
X"3a0301200093",
X"000f00000013",
X"000f00000013",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"343301f00193",
X"48c70e771263",
X"005f00000213",
X"0e3f00d00113",
X"000f00000013",
X"080300700093",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"503302000193",
X"28870a771c63",
X"005f00000213",
X"0e3f00d00113",
X"000f00000013",
X"330301300093",
X"000f00000013",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"593302100193",
X"78f708771463",
X"005f00000213",
X"0e3f00d00113",
X"000f00000013",
X"000f00000013",
X"010300600093",
X"0a650020a733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"5a3302200193",
X"688704771c63",
X"3403fff00093",
X"099500102133",
X"006300000393",
X"533302300193",
X"6bc704711263",
X"3403fff00093",
X"00550000a133",
X"096300100393",
X"5b3302400193",
X"5be702711863",
X"00a9000020b3",
X"006300000393",
X"523302500193",
X"585702709063",
X"300301000093",
X"3d3f01e00113",
X"0a650020a033",
X"006300000393",
X"513302600193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"3e66ce1fa06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6e66cc1fa06f",
X"000300000093",
X"003f00000113",
X"0af50020b733",
X"006300000393",
X"0a3300200193",
X"98b74a771a63",
X"090300100093",
X"093f00100113",
X"0af50020b733",
X"006300000393",
X"033300300193",
X"c8d748771e63",
X"030300300093",
X"083f00700113",
X"0af50020b733",
X"096300100393",
X"0b3300400193",
X"c8c748771263",
X"080300700093",
X"033f00300113",
X"0af50020b733",
X"006300000393",
X"023300500193",
X"88a746771663",
X"000300000093",
X"33f3ffff8137",
X"0af50020b733",
X"096300100393",
X"013300600193",
X"d8b744771a63",
X"c00f800000b7",
X"003f00000113",
X"0af50020b733",
X"006300000393",
X"083300700193",
X"e8d742771e63",
X"c00f800000b7",
X"33f3ffff8137",
X"0af50020b733",
X"096300100393",
X"0c3300800193",
X"e8c742771263",
X"000300000093",
X"00f300008137",
X"373ffff10113",
X"0af50020b733",
X"096300100393",
X"053300900193",
X"b8f740771463",
X"c00f800000b7",
X"34c3fff08093",
X"003f00000113",
X"0af50020b733",
X"006300000393",
X"063300a00193",
X"78a73e771663",
X"c00f800000b7",
X"34c3fff08093",
X"00f300008137",
X"373ffff10113",
X"0af50020b733",
X"006300000393",
X"0f3300b00193",
X"28a73c771663",
X"c00f800000b7",
X"00f300008137",
X"373ffff10113",
X"0af50020b733",
X"006300000393",
X"073300c00193",
X"18e73a771863",
X"c00f800000b7",
X"34c3fff08093",
X"33f3ffff8137",
X"0af50020b733",
X"096300100393",
X"0e3300d00193",
X"48b738771a63",
X"000300000093",
X"343ffff00113",
X"0af50020b733",
X"096300100393",
X"0d3300e00193",
X"08d736771e63",
X"3403fff00093",
X"093f00100113",
X"0af50020b733",
X"006300000393",
X"043300f00193",
X"08c736771263",
X"3403fff00093",
X"343ffff00113",
X"0af50020b733",
X"006300000393",
X"303301000193",
X"58a734771663",
X"0d0300e00093",
X"0e3f00d00113",
X"0af90020b0b3",
X"006300000393",
X"393301100193",
X"687732709a63",
X"0f0300b00093",
X"0e3f00d00113",
X"0ac50020b133",
X"096300100393",
X"3a3301200193",
X"3bd730711e63",
X"0e0300d00093",
X"09f90010b0b3",
X"006300000393",
X"333301300193",
X"383730709463",
X"005f00000213",
X"0f0300b00093",
X"0e3f00d00113",
X"0af50020b733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"3b3301400193",
X"bed72c731e63",
X"005f00000213",
X"0d0300e00093",
X"0e3f00d00113",
X"0af50020b733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"323301500193",
X"8ea72a731663",
X"005f00000213",
X"070300c00093",
X"0e3f00d00113",
X"0af50020b733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"096300100393",
X"313301600193",
X"9e8726731c63",
X"005f00000213",
X"0d0300e00093",
X"0e3f00d00113",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"383301700193",
X"c8e724771863",
X"005f00000213",
X"0f0300b00093",
X"0e3f00d00113",
X"000f00000013",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"3c3301800193",
X"f8c722771263",
X"005f00000213",
X"040300f00093",
X"0e3f00d00113",
X"000f00000013",
X"000f00000013",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"353301900193",
X"d8b71e771a63",
X"005f00000213",
X"060300a00093",
X"000f00000013",
X"0e3f00d00113",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"363301a00193",
X"88f71c771463",
X"005f00000213",
X"300301000093",
X"000f00000013",
X"0e3f00d00113",
X"000f00000013",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"3f3301b00193",
X"e88718771c63",
X"005f00000213",
X"050300900093",
X"000f00000013",
X"000f00000013",
X"0e3f00d00113",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"373301c00193",
X"a8f716771463",
X"005f00000213",
X"0e3f00d00113",
X"390301100093",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"006300000393",
X"3e3301d00193",
X"f89714771063",
X"005f00000213",
X"0e3f00d00113",
X"0c0300800093",
X"000f00000013",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"3d3301e00193",
X"98b710771a63",
X"005f00000213",
X"0e3f00d00113",
X"3a0301200093",
X"000f00000013",
X"000f00000013",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"343301f00193",
X"48c70e771263",
X"005f00000213",
X"0e3f00d00113",
X"000f00000013",
X"080300700093",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"096300100393",
X"503302000193",
X"28870a771c63",
X"005f00000213",
X"0e3f00d00113",
X"000f00000013",
X"330301300093",
X"000f00000013",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"006300000393",
X"593302100193",
X"78f708771463",
X"005f00000213",
X"0e3f00d00113",
X"000f00000013",
X"000f00000013",
X"010300600093",
X"0af50020b733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"5a3302200193",
X"688704771c63",
X"3403fff00093",
X"090500103133",
X"096300100393",
X"533302300193",
X"6bc704711263",
X"3403fff00093",
X"00c50000b133",
X"006300000393",
X"5b3302400193",
X"5be702711863",
X"0039000030b3",
X"006300000393",
X"523302500193",
X"585702709063",
X"300301000093",
X"3d3f01e00113",
X"0af50020b033",
X"006300000393",
X"513302600193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6066fdcfa06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"5066fbcfa06f",
X"000300000093",
X"b0ef4000d713",
X"006300000393",
X"0a3300200193",
X"88f72a771463",
X"c00f800000b7",
X"b9ef4010d713",
X"706fc00003b7",
X"033300300193",
X"d8b728771a63",
X"c00f800000b7",
X"b8ef4070d713",
X"306fff0003b7",
X"0b3300400193",
X"d89728771063",
X"c00f800000b7",
X"bdef40e0d713",
X"306ffffe03b7",
X"023300500193",
X"98a726771663",
X"c00f800000b7",
X"09c300108093",
X"84ef41f0d713",
X"3463fff00393",
X"013300600193",
X"c8b724771a63",
X"c00f800000b7",
X"34c3fff08093",
X"b0ef4000d713",
X"c06f800003b7",
X"32a3fff38393",
X"083300700193",
X"f88722771c63",
X"c00f800000b7",
X"34c3fff08093",
X"b9ef4010d713",
X"b06f400003b7",
X"32a3fff38393",
X"0c3300800193",
X"a8d720771e63",
X"c00f800000b7",
X"34c3fff08093",
X"b8ef4070d713",
X"306f010003b7",
X"32a3fff38393",
X"053300900193",
X"a89720771063",
X"c00f800000b7",
X"34c3fff08093",
X"bdef40e0d713",
X"056f000203b7",
X"32a3fff38393",
X"063300a00193",
X"d8c71e771263",
X"c00f800000b7",
X"34c3fff08093",
X"84ef41f0d713",
X"006300000393",
X"0f3300b00193",
X"88a71c771663",
X"ffcf818180b7",
X"e9c318108093",
X"b0ef4000d713",
X"ffaf818183b7",
X"efa318138393",
X"073300c00193",
X"b8e71a771863",
X"ffcf818180b7",
X"e9c318108093",
X"b9ef4010d713",
X"771fc0c0c3b7",
X"16a30c038393",
X"0e3300d00193",
X"e8b718771a63",
X"ffcf818180b7",
X"e9c318108093",
X"b8ef4070d713",
X"366fff0303b7",
X"35a330338393",
X"0d3300e00193",
X"a88716771c63",
X"ffcf818180b7",
X"e9c318108093",
X"bdef40e0d713",
X"306ffffe03b7",
X"17a360638393",
X"043300f00193",
X"f8d714771e63",
X"ffcf818180b7",
X"e9c318108093",
X"84ef41f0d713",
X"3463fff00393",
X"303301000193",
X"f8c714771263",
X"c00f800000b7",
X"b8e34070d093",
X"306fff0003b7",
X"393301100193",
X"c82712709863",
X"005f00000213",
X"c00f800000b7",
X"b8ef4070d713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306fff0003b7",
X"3a3301200193",
X"9ef710731463",
X"005f00000213",
X"c00f800000b7",
X"bdef40e0d713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306ffffe03b7",
X"333301300193",
X"1ed70c731e63",
X"005f00000213",
X"c00f800000b7",
X"09c300108093",
X"84ef41f0d713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"3463fff00393",
X"3b3301400193",
X"2ef70a731463",
X"005f00000213",
X"c00f800000b7",
X"b8ef4070d713",
X"0c5f00120213",
X"0a5300200293",
X"07ebfe5218e3",
X"306fff0003b7",
X"323301500193",
X"78c708771263",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"bdef40e0d713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306ffffe03b7",
X"313301600193",
X"68d704771e63",
X"005f00000213",
X"c00f800000b7",
X"09c300108093",
X"000f00000013",
X"000f00000013",
X"84ef41f0d713",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3463fff00393",
X"383301700193",
X"58a702771663",
X"bb2340405093",
X"006300000393",
X"3c3301800193",
X"081700709e63",
X"590302100093",
X"b6ef40a0d013",
X"006300000393",
X"353301900193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"3b66ce8fa06f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"6b66cc8fa06f",
X"c00f800000b7",
X"003f00000113",
X"bae54020d733",
X"c06f800003b7",
X"0a3300200193",
X"58f758771463",
X"c00f800000b7",
X"093f00100113",
X"bae54020d733",
X"706fc00003b7",
X"033300300193",
X"18e756771863",
X"c00f800000b7",
X"083f00700113",
X"bae54020d733",
X"306fff0003b7",
X"0b3300400193",
X"488754771c63",
X"c00f800000b7",
X"0d3f00e00113",
X"bae54020d733",
X"306ffffe03b7",
X"023300500193",
X"489754771063",
X"c00f800000b7",
X"09c300108093",
X"343f01f00113",
X"bae54020d733",
X"3463fff00393",
X"013300600193",
X"78c752771263",
X"c00f800000b7",
X"34c3fff08093",
X"003f00000113",
X"bae54020d733",
X"c06f800003b7",
X"32a3fff38393",
X"083300700193",
X"28c750771263",
X"c00f800000b7",
X"34c3fff08093",
X"093f00100113",
X"bae54020d733",
X"b06f400003b7",
X"32a3fff38393",
X"0c3300800193",
X"f8c74e771263",
X"c00f800000b7",
X"34c3fff08093",
X"083f00700113",
X"bae54020d733",
X"306f010003b7",
X"32a3fff38393",
X"053300900193",
X"a8c74c771263",
X"c00f800000b7",
X"34c3fff08093",
X"0d3f00e00113",
X"bae54020d733",
X"056f000203b7",
X"32a3fff38393",
X"063300a00193",
X"98c74a771263",
X"c00f800000b7",
X"34c3fff08093",
X"343f01f00113",
X"bae54020d733",
X"006300000393",
X"0f3300b00193",
X"c8f748771463",
X"ffcf818180b7",
X"e9c318108093",
X"003f00000113",
X"bae54020d733",
X"ffaf818183b7",
X"efa318138393",
X"073300c00193",
X"88f746771463",
X"ffcf818180b7",
X"e9c318108093",
X"093f00100113",
X"bae54020d733",
X"771fc0c0c3b7",
X"16a30c038393",
X"0e3300d00193",
X"d8f744771463",
X"ffcf818180b7",
X"e9c318108093",
X"083f00700113",
X"bae54020d733",
X"366fff0303b7",
X"35a330338393",
X"0d3300e00193",
X"e8f742771463",
X"ffcf818180b7",
X"e9c318108093",
X"0d3f00e00113",
X"bae54020d733",
X"306ffffe03b7",
X"17a360638393",
X"043300f00193",
X"b8f740771463",
X"ffcf818180b7",
X"e9c318108093",
X"343f01f00113",
X"bae54020d733",
X"3463fff00393",
X"303301000193",
X"78a73e771663",
X"ffcf818180b7",
X"e9c318108093",
X"503ffc000113",
X"bae54020d733",
X"ffaf818183b7",
X"efa318138393",
X"393301100193",
X"28a73c771663",
X"ffcf818180b7",
X"e9c318108093",
X"593ffc100113",
X"bae54020d733",
X"771fc0c0c3b7",
X"16a30c038393",
X"3a3301200193",
X"18a73a771663",
X"ffcf818180b7",
X"e9c318108093",
X"583ffc700113",
X"bae54020d733",
X"366fff0303b7",
X"35a330338393",
X"333301300193",
X"48a738771663",
X"ffcf818180b7",
X"e9c318108093",
X"5d3ffce00113",
X"bae54020d733",
X"306ffffe03b7",
X"17a360638393",
X"3b3301400193",
X"08a736771663",
X"ffcf818180b7",
X"e9c318108093",
X"343ffff00113",
X"bae54020d733",
X"3463fff00393",
X"323301500193",
X"58e734771863",
X"c00f800000b7",
X"083f00700113",
X"bae94020d0b3",
X"306fff0003b7",
X"313301600193",
X"684732709c63",
X"c00f800000b7",
X"0d3f00e00113",
X"bad54020d133",
X"306ffffe03b7",
X"383301700193",
X"6b9732711063",
X"080300700093",
X"b9e94010d0b3",
X"006300000393",
X"3c3301800193",
X"386730709663",
X"005f00000213",
X"c00f800000b7",
X"083f00700113",
X"bae54020d733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306fff0003b7",
X"353301900193",
X"ee972e731063",
X"005f00000213",
X"c00f800000b7",
X"0d3f00e00113",
X"bae54020d733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"306ffffe03b7",
X"363301a00193",
X"8ee72a731863",
X"005f00000213",
X"c00f800000b7",
X"343f01f00113",
X"bae54020d733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"3463fff00393",
X"3f3301b00193",
X"9ed726731e63",
X"005f00000213",
X"c00f800000b7",
X"083f00700113",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306fff0003b7",
X"373301c00193",
X"c8b724771a63",
X"005f00000213",
X"c00f800000b7",
X"0d3f00e00113",
X"000f00000013",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306ffffe03b7",
X"3e3301d00193",
X"f8f722771463",
X"005f00000213",
X"c00f800000b7",
X"343f01f00113",
X"000f00000013",
X"000f00000013",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3463fff00393",
X"3d3301e00193",
X"d8871e771c63",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"083f00700113",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306fff0003b7",
X"343301f00193",
X"88a71c771663",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"0d3f00e00113",
X"000f00000013",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"306ffffe03b7",
X"503302000193",
X"e8d718771e63",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"000f00000013",
X"343f01f00113",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3463fff00393",
X"593302100193",
X"a8a716771663",
X"005f00000213",
X"083f00700113",
X"c00f800000b7",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306fff0003b7",
X"5a3302200193",
X"f8c714771263",
X"005f00000213",
X"0d3f00e00113",
X"c00f800000b7",
X"000f00000013",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306ffffe03b7",
X"533302300193",
X"988710771c63",
X"005f00000213",
X"343f01f00113",
X"c00f800000b7",
X"000f00000013",
X"000f00000013",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3463fff00393",
X"5b3302400193",
X"48f70e771463",
X"005f00000213",
X"083f00700113",
X"000f00000013",
X"c00f800000b7",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306fff0003b7",
X"523302500193",
X"28d70a771e63",
X"005f00000213",
X"0d3f00e00113",
X"000f00000013",
X"c00f800000b7",
X"000f00000013",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"306ffffe03b7",
X"513302600193",
X"78a708771663",
X"005f00000213",
X"343f01f00113",
X"000f00000013",
X"000f00000013",
X"c00f800000b7",
X"bae54020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"3463fff00393",
X"583302700193",
X"68d704771e63",
X"040300f00093",
X"b91540105133",
X"006300000393",
X"5c3302800193",
X"6bf704711463",
X"500302000093",
X"b0d54000d133",
X"506302000393",
X"553302900193",
X"5bb702711a63",
X"b029400050b3",
X"006300000393",
X"563302a00193",
X"580702709263",
X"b00340000093",
X"00a300001137",
X"c33f80010113",
X"bae54020d033",
X"006300000393",
X"5f3302b00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"7e56f11f906f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"ae56ef1f906f",
X"c00f800000b7",
X"00ef0000d713",
X"c06f800003b7",
X"0a3300200193",
X"d8e728771863",
X"c00f800000b7",
X"09ef0010d713",
X"b06f400003b7",
X"033300300193",
X"98d726771e63",
X"c00f800000b7",
X"08ef0070d713",
X"306f010003b7",
X"0b3300400193",
X"98f726771463",
X"c00f800000b7",
X"0def00e0d713",
X"056f000203b7",
X"023300500193",
X"c8b724771a63",
X"c00f800000b7",
X"09c300108093",
X"34ef01f0d713",
X"096300100393",
X"013300600193",
X"f8d722771e63",
X"3403fff00093",
X"00ef0000d713",
X"3463fff00393",
X"083300700193",
X"f8f722771463",
X"3403fff00093",
X"09ef0010d713",
X"c06f800003b7",
X"32a3fff38393",
X"0c3300800193",
X"a8e720771863",
X"3403fff00093",
X"08ef0070d713",
X"506f020003b7",
X"32a3fff38393",
X"053300900193",
X"d8871e771c63",
X"3403fff00093",
X"0def00e0d713",
X"066f000403b7",
X"32a3fff38393",
X"063300a00193",
X"d8971e771063",
X"3403fff00093",
X"34ef01f0d713",
X"096300100393",
X"0f3300b00193",
X"88a71c771663",
X"99af212120b7",
X"c9c312108093",
X"00ef0000d713",
X"99cf212123b7",
X"cfa312138393",
X"073300c00193",
X"b8e71a771863",
X"99af212120b7",
X"c9c312108093",
X"09ef0010d713",
X"953f109093b7",
X"46a309038393",
X"0e3300d00193",
X"e8b718771a63",
X"99af212120b7",
X"c9c312108093",
X"08ef0070d713",
X"0edf004243b7",
X"cca324238393",
X"0d3300e00193",
X"a88716771c63",
X"99af212120b7",
X"c9c312108093",
X"0def00e0d713",
X"00af000083b7",
X"cda348438393",
X"043300f00193",
X"f8d714771e63",
X"99af212120b7",
X"c9c312108093",
X"34ef01f0d713",
X"006300000393",
X"303301000193",
X"f8c714771263",
X"c00f800000b7",
X"08e30070d093",
X"306f010003b7",
X"393301100193",
X"c82712709863",
X"005f00000213",
X"c00f800000b7",
X"08ef0070d713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306f010003b7",
X"3a3301200193",
X"9ef710731463",
X"005f00000213",
X"c00f800000b7",
X"0def00e0d713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"056f000203b7",
X"333301300193",
X"1ed70c731e63",
X"005f00000213",
X"c00f800000b7",
X"09c300108093",
X"34ef01f0d713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"096300100393",
X"3b3301400193",
X"2ef70a731463",
X"005f00000213",
X"c00f800000b7",
X"08ef0070d713",
X"0c5f00120213",
X"0a5300200293",
X"07ebfe5218e3",
X"306f010003b7",
X"323301500193",
X"78c708771263",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"0def00e0d713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"056f000203b7",
X"313301600193",
X"68d704771e63",
X"005f00000213",
X"c00f800000b7",
X"09c300108093",
X"000f00000013",
X"000f00000013",
X"34ef01f0d713",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"383301700193",
X"58a702771663",
X"0b2300405093",
X"006300000393",
X"3c3301800193",
X"081700709e63",
X"590302100093",
X"06ef00a0d013",
X"006300000393",
X"353301900193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"1556c35f906f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"4556c15f906f",
X"c00f800000b7",
X"003f00000113",
X"0ae50020d733",
X"c06f800003b7",
X"0a3300200193",
X"18e756771863",
X"c00f800000b7",
X"093f00100113",
X"0ae50020d733",
X"b06f400003b7",
X"033300300193",
X"488754771c63",
X"c00f800000b7",
X"083f00700113",
X"0ae50020d733",
X"306f010003b7",
X"0b3300400193",
X"489754771063",
X"c00f800000b7",
X"0d3f00e00113",
X"0ae50020d733",
X"056f000203b7",
X"023300500193",
X"78f752771463",
X"c00f800000b7",
X"09c300108093",
X"343f01f00113",
X"0ae50020d733",
X"096300100393",
X"013300600193",
X"28a750771663",
X"3403fff00093",
X"003f00000113",
X"0ae50020d733",
X"3463fff00393",
X"083300700193",
X"f8b74e771a63",
X"3403fff00093",
X"093f00100113",
X"0ae50020d733",
X"c06f800003b7",
X"32a3fff38393",
X"0c3300800193",
X"a8874c771c63",
X"3403fff00093",
X"083f00700113",
X"0ae50020d733",
X"506f020003b7",
X"32a3fff38393",
X"053300900193",
X"98d74a771e63",
X"3403fff00093",
X"0d3f00e00113",
X"0ae50020d733",
X"066f000403b7",
X"32a3fff38393",
X"063300a00193",
X"98974a771063",
X"3403fff00093",
X"343f01f00113",
X"0ae50020d733",
X"096300100393",
X"0f3300b00193",
X"c8f748771463",
X"99af212120b7",
X"c9c312108093",
X"003f00000113",
X"0ae50020d733",
X"99cf212123b7",
X"cfa312138393",
X"073300c00193",
X"88f746771463",
X"99af212120b7",
X"c9c312108093",
X"093f00100113",
X"0ae50020d733",
X"953f109093b7",
X"46a309038393",
X"0e3300d00193",
X"d8f744771463",
X"99af212120b7",
X"c9c312108093",
X"083f00700113",
X"0ae50020d733",
X"0edf004243b7",
X"cca324238393",
X"0d3300e00193",
X"e8f742771463",
X"99af212120b7",
X"c9c312108093",
X"0d3f00e00113",
X"0ae50020d733",
X"00af000083b7",
X"cda348438393",
X"043300f00193",
X"b8f740771463",
X"99af212120b7",
X"c9c312108093",
X"343f01f00113",
X"0ae50020d733",
X"006300000393",
X"303301000193",
X"78a73e771663",
X"99af212120b7",
X"c9c312108093",
X"503ffc000113",
X"0ae50020d733",
X"99cf212123b7",
X"cfa312138393",
X"393301100193",
X"28a73c771663",
X"99af212120b7",
X"c9c312108093",
X"593ffc100113",
X"0ae50020d733",
X"953f109093b7",
X"46a309038393",
X"3a3301200193",
X"18a73a771663",
X"99af212120b7",
X"c9c312108093",
X"583ffc700113",
X"0ae50020d733",
X"0edf004243b7",
X"cca324238393",
X"333301300193",
X"48a738771663",
X"99af212120b7",
X"c9c312108093",
X"5d3ffce00113",
X"0ae50020d733",
X"00af000083b7",
X"cda348438393",
X"3b3301400193",
X"08a736771663",
X"99af212120b7",
X"c9c312108093",
X"343ffff00113",
X"0ae50020d733",
X"006300000393",
X"323301500193",
X"58e734771863",
X"c00f800000b7",
X"083f00700113",
X"0ae90020d0b3",
X"306f010003b7",
X"313301600193",
X"684732709c63",
X"c00f800000b7",
X"0d3f00e00113",
X"0ad50020d133",
X"056f000203b7",
X"383301700193",
X"6b9732711063",
X"080300700093",
X"09e90010d0b3",
X"006300000393",
X"3c3301800193",
X"386730709663",
X"005f00000213",
X"c00f800000b7",
X"083f00700113",
X"0ae50020d733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306f010003b7",
X"353301900193",
X"ee972e731063",
X"005f00000213",
X"c00f800000b7",
X"0d3f00e00113",
X"0ae50020d733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"056f000203b7",
X"363301a00193",
X"8ee72a731863",
X"005f00000213",
X"c00f800000b7",
X"343f01f00113",
X"0ae50020d733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"096300100393",
X"3f3301b00193",
X"9ed726731e63",
X"005f00000213",
X"c00f800000b7",
X"083f00700113",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306f010003b7",
X"373301c00193",
X"c8b724771a63",
X"005f00000213",
X"c00f800000b7",
X"0d3f00e00113",
X"000f00000013",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"056f000203b7",
X"3e3301d00193",
X"f8f722771463",
X"005f00000213",
X"c00f800000b7",
X"343f01f00113",
X"000f00000013",
X"000f00000013",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"3d3301e00193",
X"d8871e771c63",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"083f00700113",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306f010003b7",
X"343301f00193",
X"88a71c771663",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"0d3f00e00113",
X"000f00000013",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"056f000203b7",
X"503302000193",
X"e8d718771e63",
X"005f00000213",
X"c00f800000b7",
X"000f00000013",
X"000f00000013",
X"343f01f00113",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"593302100193",
X"a8a716771663",
X"005f00000213",
X"083f00700113",
X"c00f800000b7",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"306f010003b7",
X"5a3302200193",
X"f8c714771263",
X"005f00000213",
X"0d3f00e00113",
X"c00f800000b7",
X"000f00000013",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"056f000203b7",
X"533302300193",
X"988710771c63",
X"005f00000213",
X"343f01f00113",
X"c00f800000b7",
X"000f00000013",
X"000f00000013",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"5b3302400193",
X"48f70e771463",
X"005f00000213",
X"083f00700113",
X"000f00000013",
X"c00f800000b7",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"306f010003b7",
X"523302500193",
X"28d70a771e63",
X"005f00000213",
X"0d3f00e00113",
X"000f00000013",
X"c00f800000b7",
X"000f00000013",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"056f000203b7",
X"513302600193",
X"78a708771663",
X"005f00000213",
X"343f01f00113",
X"000f00000013",
X"000f00000013",
X"c00f800000b7",
X"0ae50020d733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"096300100393",
X"583302700193",
X"68d704771e63",
X"040300f00093",
X"091500105133",
X"006300000393",
X"5c3302800193",
X"6bf704711463",
X"500302000093",
X"00d50000d133",
X"506302000393",
X"553302900193",
X"5bb702711a63",
X"0029000050b3",
X"006300000393",
X"563302a00193",
X"580702709263",
X"b00340000093",
X"00a300001137",
X"c33f80010113",
X"0ae50020d033",
X"006300000393",
X"5f3302b00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"dc56e74f906f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"8c56e54f906f",
X"000300000093",
X"003f00000113",
X"bac540208733",
X"006300000393",
X"0a3300200193",
X"98a74a771663",
X"090300100093",
X"093f00100113",
X"bac540208733",
X"006300000393",
X"033300300193",
X"c8b748771a63",
X"030300300093",
X"083f00700113",
X"bac540208733",
X"3763ffc00393",
X"0b3300400193",
X"88d746771e63",
X"000300000093",
X"33f3ffff8137",
X"bac540208733",
X"00af000083b7",
X"023300500193",
X"88c746771263",
X"c00f800000b7",
X"003f00000113",
X"bac540208733",
X"c06f800003b7",
X"013300600193",
X"d8a744771663",
X"c00f800000b7",
X"33f3ffff8137",
X"bac540208733",
X"c0af800083b7",
X"083300700193",
X"e8b742771a63",
X"000300000093",
X"00f300008137",
X"373ffff10113",
X"bac540208733",
X"33afffff83b7",
X"0fa300138393",
X"0c3300800193",
X"b8b740771a63",
X"c00f800000b7",
X"34c3fff08093",
X"003f00000113",
X"bac540208733",
X"c06f800003b7",
X"32a3fff38393",
X"053300900193",
X"78b73e771a63",
X"c00f800000b7",
X"34c3fff08093",
X"00f300008137",
X"373ffff10113",
X"bac540208733",
X"f3af7fff83b7",
X"063300a00193",
X"28b73c771a63",
X"c00f800000b7",
X"00f300008137",
X"373ffff10113",
X"bac540208733",
X"f3af7fff83b7",
X"0fa300138393",
X"0f3300b00193",
X"18b73a771a63",
X"c00f800000b7",
X"34c3fff08093",
X"33f3ffff8137",
X"bac540208733",
X"c0af800083b7",
X"32a3fff38393",
X"073300c00193",
X"48b738771a63",
X"000300000093",
X"343ffff00113",
X"bac540208733",
X"096300100393",
X"0e3300d00193",
X"08d736771e63",
X"3403fff00093",
X"093f00100113",
X"bac540208733",
X"3d63ffe00393",
X"0d3300e00193",
X"08c736771263",
X"3403fff00093",
X"343ffff00113",
X"bac540208733",
X"006300000393",
X"043300f00193",
X"58a734771663",
X"0e0300d00093",
X"0f3f00b00113",
X"bac9402080b3",
X"0a6300200393",
X"303301000193",
X"687732709a63",
X"0d0300e00093",
X"0f3f00b00113",
X"baf540208133",
X"036300300393",
X"393301100193",
X"3bd730711e63",
X"0e0300d00093",
X"b9c9401080b3",
X"006300000393",
X"3a3301200193",
X"383730709463",
X"005f00000213",
X"0e0300d00093",
X"0f3f00b00113",
X"bac540208733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0a6300200393",
X"333301300193",
X"bed72c731e63",
X"005f00000213",
X"0d0300e00093",
X"0f3f00b00113",
X"bac540208733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"036300300393",
X"3b3301400193",
X"8ea72a731663",
X"005f00000213",
X"040300f00093",
X"0f3f00b00113",
X"bac540208733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"0b6300400393",
X"323301500193",
X"9e8726731c63",
X"005f00000213",
X"0e0300d00093",
X"0f3f00b00113",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"0a6300200393",
X"313301600193",
X"c8e724771863",
X"005f00000213",
X"0d0300e00093",
X"0f3f00b00113",
X"000f00000013",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"036300300393",
X"383301700193",
X"f8c722771263",
X"005f00000213",
X"040300f00093",
X"0f3f00b00113",
X"000f00000013",
X"000f00000013",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0b6300400393",
X"3c3301800193",
X"d8b71e771a63",
X"005f00000213",
X"0e0300d00093",
X"000f00000013",
X"0f3f00b00113",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0a6300200393",
X"353301900193",
X"88f71c771463",
X"005f00000213",
X"0d0300e00093",
X"000f00000013",
X"0f3f00b00113",
X"000f00000013",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"036300300393",
X"363301a00193",
X"e88718771c63",
X"005f00000213",
X"040300f00093",
X"000f00000013",
X"000f00000013",
X"0f3f00b00113",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0b6300400393",
X"3f3301b00193",
X"a8f716771463",
X"005f00000213",
X"0f3f00b00113",
X"0e0300d00093",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"0a6300200393",
X"373301c00193",
X"f89714771063",
X"005f00000213",
X"0f3f00b00113",
X"0d0300e00093",
X"000f00000013",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"036300300393",
X"3e3301d00193",
X"98b710771a63",
X"005f00000213",
X"0f3f00b00113",
X"040300f00093",
X"000f00000013",
X"000f00000013",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0b6300400393",
X"3d3301e00193",
X"48c70e771263",
X"005f00000213",
X"0f3f00b00113",
X"000f00000013",
X"0e0300d00093",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"0a6300200393",
X"343301f00193",
X"28870a771c63",
X"005f00000213",
X"0f3f00b00113",
X"000f00000013",
X"0d0300e00093",
X"000f00000013",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"036300300393",
X"503302000193",
X"78f708771463",
X"005f00000213",
X"0f3f00b00113",
X"000f00000013",
X"000f00000013",
X"040300f00093",
X"bac540208733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"0b6300400393",
X"593302100193",
X"688704771c63",
X"3903ff100093",
X"b93540100133",
X"046300f00393",
X"5a3302200193",
X"6bc704711263",
X"500302000093",
X"b0f540008133",
X"506302000393",
X"533302300193",
X"5be702711863",
X"b009400000b3",
X"006300000393",
X"5b3302400193",
X"585702709063",
X"300301000093",
X"3d3f01e00113",
X"bac540208033",
X"006300000393",
X"523302500193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"5b56978f906f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"0b56958f906f",
X"700308000093",
X"043300aa0137",
X"253f0aa10113",
X"0a6c0020a023",
X"00660000a703",
X"046f00aa03b7",
X"20a30aa38393",
X"0a3300200193",
X"b8f740771463",
X"700308000093",
X"40c3aa00b137",
X"633fa0010113",
X"0a3c0020a223",
X"0b660040a703",
X"409faa00b3b7",
X"66a3a0038393",
X"033300300193",
X"78c73e771263",
X"700308000093",
X"26a30aa01137",
X"433faa010113",
X"0a0c0020a423",
X"0c660080a703",
X"26ff0aa013b7",
X"46a3aa038393",
X"0b3300400193",
X"28973c771063",
X"700308000093",
X"6253a00aa137",
X"053f00a10113",
X"0a5c0020a623",
X"076600c0a703",
X"620fa00aa3b7",
X"00a300a38393",
X"023300500193",
X"48d738771e63",
X"470309c00093",
X"043300aa0137",
X"253f0aa10113",
X"0a4cfe20aa23",
X"3b66ff40a703",
X"046f00aa03b7",
X"20a30aa38393",
X"013300600193",
X"088736771c63",
X"470309c00093",
X"40c3aa00b137",
X"633fa0010113",
X"0a7cfe20ac23",
X"3c66ff80a703",
X"409faa00b3b7",
X"66a3a0038393",
X"083300700193",
X"58b734771a63",
X"470309c00093",
X"26a30aa01137",
X"433faa010113",
X"0a2cfe20ae23",
X"3766ffc0a703",
X"26ff0aa013b7",
X"46a3aa038393",
X"0c3300800193",
X"68e732771863",
X"470309c00093",
X"6253a00aa137",
X"053f00a10113",
X"0a6c0020a023",
X"00660000a703",
X"620fa00aa3b7",
X"00a300a38393",
X"053300900193",
X"38a730771663",
X"20030a000093",
X"c51312345137",
X"1f3f67810113",
X"009ffe008213",
X"5fac02222023",
X"003a0000a283",
X"c54f123453b7",
X"1aa367838393",
X"063300a00193",
X"ed072e729263",
X"20030a000093",
X"590358213137",
X"4f3f09810113",
X"3ec3ffd08093",
X"0a000020a3a3",
X"2b5f0a400213",
X"05fa00022283",
X"595f582133b7",
X"4aa309838393",
X"0f3300b00193",
X"8d472a729c63",
X"073300c00193",
X"005f00000213",
X"4eefaabbd0b7",
X"5ec3cdd08093",
X"703f08000113",
X"0aac00112023",
X"03a600012703",
X"4e8faabbd3b7",
X"58a3cdd38393",
X"d8e728771863",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"0e3300d00193",
X"005f00000213",
X"c77fdaabc0b7",
X"6ec3ccd08093",
X"703f08000113",
X"000f00000013",
X"0afc00112223",
X"08a600412703",
X"c71fdaabc3b7",
X"68a3ccd38393",
X"c88724771c63",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"0d3300e00193",
X"005f00000213",
X"c47fddaac0b7",
X"e7c3bcc08093",
X"703f08000113",
X"000f00000013",
X"000f00000013",
X"0acc00112423",
X"0fa600812703",
X"c41fddaac3b7",
X"e1a3bcc38393",
X"a8d720771e63",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"043300f00193",
X"005f00000213",
X"5cffcddab0b7",
X"e7c3bbc08093",
X"000f00000013",
X"703f08000113",
X"0a9c00112623",
X"04a600c12703",
X"5c9fcddab3b7",
X"e1a3bbc38393",
X"d8c71e771263",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"303301000193",
X"005f00000213",
X"6cffccddb0b7",
X"7fc3abb08093",
X"000f00000013",
X"703f08000113",
X"000f00000013",
X"0adc00112823",
X"33a601012703",
X"6c9fccddb3b7",
X"79a3abb38393",
X"b8f71a771463",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"393301100193",
X"005f00000213",
X"e5dfbccde0b7",
X"4fc3aab08093",
X"000f00000013",
X"000f00000013",
X"703f08000113",
X"0a8c00112a23",
X"38a601412703",
X"e5bfbccde3b7",
X"49a3aab38393",
X"a8a716771663",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"3a3301200193",
X"005f00000213",
X"703f08000113",
X"0aaf001120b7",
X"c3c323308093",
X"0aac00112023",
X"03a600012703",
X"0acf001123b7",
X"c5a323338393",
X"c88712771c63",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"333301300193",
X"005f00000213",
X"703f08000113",
X"339f300110b7",
X"f3c322308093",
X"000f00000013",
X"0afc00112223",
X"08a600412703",
X"33ff300113b7",
X"f5a322338393",
X"989710771063",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"3b3301400193",
X"005f00000213",
X"703f08000113",
X"509f330010b7",
X"cac312208093",
X"000f00000013",
X"000f00000013",
X"0acc00112423",
X"0fa600812703",
X"50ff330013b7",
X"cca312238393",
X"18c70c771263",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"323301500193",
X"005f00000213",
X"703f08000113",
X"000f00000013",
X"c30f233000b7",
X"aac311208093",
X"0a9c00112623",
X"04a600c12703",
X"c36f233003b7",
X"aca311238393",
X"78a708771663",
X"0c5f00120213",
X"0a5300200293",
X"57bbfc521ae3",
X"313301600193",
X"005f00000213",
X"703f08000113",
X"000f00000013",
X"f50f223300b7",
X"39c301108093",
X"000f00000013",
X"0adc00112823",
X"33a601012703",
X"f56f223303b7",
X"3fa301138393",
X"68e704771863",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"383301700193",
X"005f00000213",
X"703f08000113",
X"000f00000013",
X"000f00000013",
X"cc3f122330b7",
X"09c300108093",
X"0a8c00112a23",
X"38a601412703",
X"cc5f122333b7",
X"0fa300138393",
X"08b700771a63",
X"0c5f00120213",
X"0a5300200293",
X"57ebfc5218e3",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"d5c6d15f806f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"05c6cf5f806f",
X"039f00ff10b7",
X"40c3f0008093",
X"447ff0f0c713",
X"302fff00f3b7",
X"02a300f38393",
X"0a3300200193",
X"88a71c771663",
X"749f0ff010b7",
X"30c3ff008093",
X"707f0f00c713",
X"74ff0ff013b7",
X"46a3f0038393",
X"033300300193",
X"b8e71a771863",
X"039f00ff10b7",
X"b4c38ff08093",
X"847f70f0c713",
X"03ff00ff13b7",
X"36a3ff038393",
X"0b3300400193",
X"e8b718771a63",
X"474ff00ff0b7",
X"04c300f08093",
X"707f0f00c713",
X"472ff00ff3b7",
X"72a30ff38393",
X"023300500193",
X"a88716771c63",
X"304fff00f0b7",
X"80c370008093",
X"847370f0c093",
X"302fff00f3b7",
X"02a300f38393",
X"013300600193",
X"f81714709e63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"707f0f00c713",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"74ff0ff013b7",
X"46a3f0038393",
X"083300700193",
X"cea712731663",
X"005f00000213",
X"039f00ff10b7",
X"b4c38ff08093",
X"847f70f0c713",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"03ff00ff13b7",
X"36a3ff038393",
X"0c3300800193",
X"4e870e731c63",
X"005f00000213",
X"474ff00ff0b7",
X"04c300f08093",
X"707f0f00c713",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"472ff00ff3b7",
X"72a30ff38393",
X"053300900193",
X"1e970c731063",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"707f0f00c713",
X"0c5f00120213",
X"0a5300200293",
X"07abfe5216e3",
X"74ff0ff013b7",
X"46a3f0038393",
X"063300a00193",
X"78b708771a63",
X"005f00000213",
X"039f00ff10b7",
X"34c3fff08093",
X"000f00000013",
X"047f00f0c713",
X"0c5f00120213",
X"0a5300200293",
X"07fbfe5214e3",
X"03ff00ff13b7",
X"36a3ff038393",
X"0f3300b00193",
X"38c706771263",
X"005f00000213",
X"474ff00ff0b7",
X"04c300f08093",
X"000f00000013",
X"000f00000013",
X"707f0f00c713",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"472ff00ff3b7",
X"72a30ff38393",
X"073300c00193",
X"58e702771863",
X"70b30f004093",
X"70630f000393",
X"0e3300d00193",
X"585702709063",
X"030f00ff00b7",
X"74c30ff08093",
X"847f70f0c013",
X"006300000393",
X"0d3300e00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"15c6af5f806f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"45c6ad5f806f",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"472ff00ff3b7",
X"02a300f38393",
X"0a3300200193",
X"98974a771063",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0a750020c733",
X"336fff0103b7",
X"46a3f0038393",
X"033300300193",
X"88d746771e63",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"74ff0ff013b7",
X"36a3ff038393",
X"0b3300400193",
X"d88744771c63",
X"474ff00ff0b7",
X"04c300f08093",
X"4473f0f0f137",
X"733f0f010113",
X"0a750020c733",
X"036f00ff03b7",
X"72a30ff38393",
X"023300500193",
X"e8b742771a63",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a790020c0b3",
X"472ff00ff3b7",
X"02a300f38393",
X"013300600193",
X"b82740709863",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a450020c133",
X"472ff00ff3b7",
X"02a300f38393",
X"083300700193",
X"7ba73e711663",
X"330fff0100b7",
X"40c3f0008093",
X"09790010c0b3",
X"006300000393",
X"0c3300800193",
X"28773c709a63",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"472ff00ff3b7",
X"02a300f38393",
X"053300900193",
X"4ed738731e63",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"0a750020c733",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"336fff0103b7",
X"46a3f0038393",
X"063300a00193",
X"0e9736731063",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"000f00000013",
X"000f00000013",
X"006f00070313",
X"0c5f00120213",
X"0a5300200293",
X"578bfc521ce3",
X"74ff0ff013b7",
X"36a3ff038393",
X"0f3300b00193",
X"6e9732731063",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"472ff00ff3b7",
X"02a300f38393",
X"073300c00193",
X"e8a72e771663",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"336fff0103b7",
X"46a3f0038393",
X"0e3300d00193",
X"88b72a771a63",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"000f00000013",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"74ff0ff013b7",
X"36a3ff038393",
X"0d3300e00193",
X"988726771c63",
X"005f00000213",
X"330fff0100b7",
X"40c3f0008093",
X"000f00000013",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"472ff00ff3b7",
X"02a300f38393",
X"043300f00193",
X"c89724771063",
X"005f00000213",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"336fff0103b7",
X"46a3f0038393",
X"303301000193",
X"a8c720771263",
X"005f00000213",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"000f00000013",
X"77a30f0f1137",
X"473ff0f10113",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"74ff0ff013b7",
X"36a3ff038393",
X"393301100193",
X"88f71c771463",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"330fff0100b7",
X"40c3f0008093",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"07cbfe5212e3",
X"472ff00ff3b7",
X"02a300f38393",
X"3a3301200193",
X"e8b718771a63",
X"005f00000213",
X"4473f0f0f137",
X"733f0f010113",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"336fff0103b7",
X"46a3f0038393",
X"333301300193",
X"f8d714771e63",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"030f00ff00b7",
X"74c30ff08093",
X"000f00000013",
X"000f00000013",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"74ff0ff013b7",
X"36a3ff038393",
X"3b3301400193",
X"c89712771063",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"330fff0100b7",
X"40c3f0008093",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"079bfe5210e3",
X"472ff00ff3b7",
X"02a300f38393",
X"323301500193",
X"48f70e771463",
X"005f00000213",
X"4473f0f0f137",
X"733f0f010113",
X"000f00000013",
X"749f0ff010b7",
X"30c3ff008093",
X"000f00000013",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"336fff0103b7",
X"46a3f0038393",
X"313301600193",
X"28a70a771663",
X"005f00000213",
X"77a30f0f1137",
X"473ff0f10113",
X"000f00000013",
X"000f00000013",
X"030f00ff00b7",
X"74c30ff08093",
X"0a750020c733",
X"0c5f00120213",
X"0a5300200293",
X"57dbfc521ee3",
X"74ff0ff013b7",
X"36a3ff038393",
X"383301700193",
X"38e706771863",
X"330fff0100b7",
X"40c3f0008093",
X"098500104133",
X"336fff0103b7",
X"46a3f0038393",
X"3c3301800193",
X"6bb704711a63",
X"030f00ff00b7",
X"74c30ff08093",
X"00450000c133",
X"036f00ff03b7",
X"72a30ff38393",
X"353301900193",
X"5b8702711c63",
X"00b9000040b3",
X"006300000393",
X"363301a00193",
X"583702709463",
X"aa9f111110b7",
X"a9c311108093",
X"ff9322222137",
X"f93f22210113",
X"0a750020c033",
X"006300000393",
X"3f3301b00193",
X"08f700701463",
X"53c702301263",
X"039f00018513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"9bc6df8f806f",
X"005f00000513",
X"00ff000022b7",
X"059300028293",
X"05060002a303",
X"00ac00a32023",
X"0d6f00430313",
X"046c0062a023",
X"cbc6dd8f806f",
others => X"000000000000"
);

begin

process(clka)
begin
    if(clka'event and clka = '1') then
        if(ena = '1') then
            for i in 0 to C_NB_COL-1 loop
                if wea(i) = '1' then
                    ram_name(to_integer(unsigned(addra)))((i+1)*C_COL_WIDTH-1 downto i*C_COL_WIDTH) <= dina((i+1)*C_COL_WIDTH-1 downto i*C_COL_WIDTH);
                end if;
            end loop;
            ram_data <= ram_name(to_integer(unsigned(addra)));
        end if;
    end if;
end process;

douta <= ram_data;
 
end rtl;

