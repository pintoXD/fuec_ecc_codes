/* verilator lint_off DECLFILENAME */
module syndrome_to_flip_mask_48_16 (
    input  wire [15:0] syndrome_bin,
    output reg  [47:0] flip_mask_bin
);
    always @* begin
        case (syndrome_bin)
            16'b0000000000000001: flip_mask_bin = 48'b000000000000000100000000000000000000000000000000; // 1
            16'b0000000000000010: flip_mask_bin = 48'b000000000000001000000000000000000000000000000000; // 2
            16'b0000000000000011: flip_mask_bin = 48'b000000000000001100000000000000000000000000000000; // 3
            16'b0000000000000100: flip_mask_bin = 48'b000000000000010000000000000000000000000000000000; // 4
            16'b0000000000000101: flip_mask_bin = 48'b000000000000010100000000000000000000000000000000; // 5
            16'b0000000000000110: flip_mask_bin = 48'b000000000000011000000000000000000000000000000000; // 6
            16'b0000000000000111: flip_mask_bin = 48'b000000000000011100000000000000000000000000000000; // 7
            16'b0000000000001000: flip_mask_bin = 48'b000000000000100000000000000000000000000000000000; // 8
            16'b0000000000001001: flip_mask_bin = 48'b000000000000100100000000000000000000000000000000; // 9
            16'b0000000000001010: flip_mask_bin = 48'b000000000000101000000000000000000000000000000000; // 10
            16'b0000000000001011: flip_mask_bin = 48'b000000000000101100000000000000000000000000000000; // 11
            16'b0000000000001100: flip_mask_bin = 48'b000000000000110000000000000000000000000000000000; // 12
            16'b0000000000001101: flip_mask_bin = 48'b000000000000110100000000000000000000000000000000; // 13
            16'b0000000000001110: flip_mask_bin = 48'b000000000000111000000000000000000000000000000000; // 14
            16'b0000000000001111: flip_mask_bin = 48'b000000000000111100000000000000000000000000000000; // 15
            16'b0000000000010000: flip_mask_bin = 48'b000000000001000000000000000000000000000000000000; // 16
            16'b0000000000010010: flip_mask_bin = 48'b000000000001001000000000000000000000000000000000; // 18
            16'b0000000000010100: flip_mask_bin = 48'b000000000001010000000000000000000000000000000000; // 20
            16'b0000000000010110: flip_mask_bin = 48'b000000000001011000000000000000000000000000000000; // 22
            16'b0000000000011000: flip_mask_bin = 48'b000000000001100000000000000000000000000000000000; // 24
            16'b0000000000011010: flip_mask_bin = 48'b000000000001101000000000000000000000000000000000; // 26
            16'b0000000000011100: flip_mask_bin = 48'b000000000001110000000000000000000000000000000000; // 28
            16'b0000000000011110: flip_mask_bin = 48'b000000000001111000000000000000000000000000000000; // 30
            16'b0000000000100000: flip_mask_bin = 48'b000000000010000000000000000000000000000000000000; // 32
            16'b0000000000100100: flip_mask_bin = 48'b000000000010010000000000000000000000000000000000; // 36
            16'b0000000000101000: flip_mask_bin = 48'b000000000010100000000000000000000000000000000000; // 40
            16'b0000000000101100: flip_mask_bin = 48'b000000000010110000000000000000000000000000000000; // 44
            16'b0000000000110000: flip_mask_bin = 48'b000000000011000000000000000000000000000000000000; // 48
            16'b0000000000110100: flip_mask_bin = 48'b000000000011010000000000000000000000000000000000; // 52
            16'b0000000000111000: flip_mask_bin = 48'b000000000011100000000000000000000000000000000000; // 56
            16'b0000000000111100: flip_mask_bin = 48'b000000000011110000000000000000000000000000000000; // 60
            16'b0000000001000000: flip_mask_bin = 48'b000000000100000000000000000000000000000000000000; // 64
            16'b0000000001001000: flip_mask_bin = 48'b000000000100100000000000000000000000000000000000; // 72
            16'b0000000001010000: flip_mask_bin = 48'b000000000101000000000000000000000000000000000000; // 80
            16'b0000000001011000: flip_mask_bin = 48'b000000000101100000000000000000000000000000000000; // 88
            16'b0000000001100000: flip_mask_bin = 48'b000000000110000000000000000000000000000000000000; // 96
            16'b0000000001101000: flip_mask_bin = 48'b000000000110100000000000000000000000000000000000; // 104
            16'b0000000001110000: flip_mask_bin = 48'b000000000111000000000000000000000000000000000000; // 112
            16'b0000000001111000: flip_mask_bin = 48'b000000000111100000000000000000000000000000000000; // 120
            16'b0000000010000000: flip_mask_bin = 48'b000000001000000000000000000000000000000000000000; // 128
            16'b0000000010010000: flip_mask_bin = 48'b000000001001000000000000000000000000000000000000; // 144
            16'b0000000010100000: flip_mask_bin = 48'b000000001010000000000000000000000000000000000000; // 160
            16'b0000000010110000: flip_mask_bin = 48'b000000001011000000000000000000000000000000000000; // 176
            16'b0000000011000000: flip_mask_bin = 48'b000000001100000000000000000000000000000000000000; // 192
            16'b0000000011010000: flip_mask_bin = 48'b000000001101000000000000000000000000000000000000; // 208
            16'b0000000011100000: flip_mask_bin = 48'b000000001110000000000000000000000000000000000000; // 224
            16'b0000000011110000: flip_mask_bin = 48'b000000001111000000000000000000000000000000000000; // 240
            16'b0000000100000000: flip_mask_bin = 48'b000000010000000000000000000000000000000000000000; // 256
            16'b0000000100100000: flip_mask_bin = 48'b000000010010000000000000000000000000000000000000; // 288
            16'b0000000100111101: flip_mask_bin = 48'b000000000000000000000000000001000000000000000000; // 317
            16'b0000000101000000: flip_mask_bin = 48'b000000010100000000000000000000000000000000000000; // 320
            16'b0000000101100000: flip_mask_bin = 48'b000000010110000000000000000000000000000000000000; // 352
            16'b0000000110000000: flip_mask_bin = 48'b000000011000000000000000000000000000000000000000; // 384
            16'b0000000110100000: flip_mask_bin = 48'b000000011010000000000000000000000000000000000000; // 416
            16'b0000000111000000: flip_mask_bin = 48'b000000011100000000000000000000000000000000000000; // 448
            16'b0000000111100000: flip_mask_bin = 48'b000000011110000000000000000000000000000000000000; // 480
            16'b0000000111101010: flip_mask_bin = 48'b000000000000000000000000000000001010000000000000; // 490
            16'b0000001000000000: flip_mask_bin = 48'b000000100000000000000000000000000000000000000000; // 512
            16'b0000001001000000: flip_mask_bin = 48'b000000100100000000000000000000000000000000000000; // 576
            16'b0000001010000000: flip_mask_bin = 48'b000000101000000000000000000000000000000000000000; // 640
            16'b0000001011000000: flip_mask_bin = 48'b000000101100000000000000000000000000000000000000; // 704
            16'b0000001100000000: flip_mask_bin = 48'b000000110000000000000000000000000000000000000000; // 768
            16'b0000001100011011: flip_mask_bin = 48'b000000000000000000000001110000000000000000000000; // 795
            16'b0000001101000000: flip_mask_bin = 48'b000000110100000000000000000000000000000000000000; // 832
            16'b0000001110000000: flip_mask_bin = 48'b000000111000000000000000000000000000000000000000; // 896
            16'b0000001111000000: flip_mask_bin = 48'b000000111100000000000000000000000000000000000000; // 960
            16'b0000010000000000: flip_mask_bin = 48'b000001000000000000000000000000000000000000000000; // 1024
            16'b0000010000000111: flip_mask_bin = 48'b000000000000000000000000000000000000000010010000; // 1031
            16'b0000010010000000: flip_mask_bin = 48'b000001001000000000000000000000000000000000000000; // 1152
            16'b0000010100000000: flip_mask_bin = 48'b000001010000000000000000000000000000000000000000; // 1280
            16'b0000010110000000: flip_mask_bin = 48'b000001011000000000000000000000000000000000000000; // 1408
            16'b0000011000000000: flip_mask_bin = 48'b000001100000000000000000000000000000000000000000; // 1536
            16'b0000011001010001: flip_mask_bin = 48'b000000000000000000000000000000000000000000101100; // 1617
            16'b0000011010000000: flip_mask_bin = 48'b000001101000000000000000000000000000000000000000; // 1664
            16'b0000011010011000: flip_mask_bin = 48'b000000000000000000000000000000000000000000000001; // 1688
            16'b0000011011101000: flip_mask_bin = 48'b000000000000000000000000000000000000000110100000; // 1768
            16'b0000011100000000: flip_mask_bin = 48'b000001110000000000000000000000000000000000000000; // 1792
            16'b0000011110000000: flip_mask_bin = 48'b000001111000000000000000000000000000000000000000; // 1920
            16'b0000100000000000: flip_mask_bin = 48'b000010000000000000000000000000000000000000000000; // 2048
            16'b0000100100000000: flip_mask_bin = 48'b000010010000000000000000000000000000000000000000; // 2304
            16'b0000100101100101: flip_mask_bin = 48'b000000000000000000000000000000000000000000000111; // 2405
            16'b0000101000000000: flip_mask_bin = 48'b000010100000000000000000000000000000000000000000; // 2560
            16'b0000101001100010: flip_mask_bin = 48'b000000000000000000001000000000000000000000000000; // 2658
            16'b0000101100000000: flip_mask_bin = 48'b000010110000000000000000000000000000000000000000; // 2816
            16'b0000101110101001: flip_mask_bin = 48'b000000000000000000000000000000000000001011000000; // 2985
            16'b0000110000000000: flip_mask_bin = 48'b000011000000000000000000000000000000000000000000; // 3072
            16'b0000110100000000: flip_mask_bin = 48'b000011010000000000000000000000000000000000000000; // 3328
            16'b0000111000000000: flip_mask_bin = 48'b000011100000000000000000000000000000000000000000; // 3584
            16'b0000111100000000: flip_mask_bin = 48'b000011110000000000000000000000000000000000000000; // 3840
            16'b0000111111111101: flip_mask_bin = 48'b000000000000000000000000000000000000000000000110; // 4093
            16'b0001000000000000: flip_mask_bin = 48'b000100000000000000000000000000000000000000000000; // 4096
            16'b0001000001011110: flip_mask_bin = 48'b000000000000000000000000000000000000000001000000; // 4190
            16'b0001001000000000: flip_mask_bin = 48'b000100100000000000000000000000000000000000000000; // 4608
            16'b0001010000000000: flip_mask_bin = 48'b000101000000000000000000000000000000000000000000; // 5120
            16'b0001010000000001: flip_mask_bin = 48'b000000000000000000000000100100000000000000000000; // 5121
            16'b0001010001011001: flip_mask_bin = 48'b000000000000000000000000000000000000000011010000; // 5209
            16'b0001011000000000: flip_mask_bin = 48'b000101100000000000000000000000000000000000000000; // 5632
            16'b0001011000111110: flip_mask_bin = 48'b000000000000000000000000000001001000000000000000; // 5694
            16'b0001011010110110: flip_mask_bin = 48'b000000000000000000000000000000000000000111100000; // 5814
            16'b0001011011101001: flip_mask_bin = 48'b000000000000000000000000000000000010000000000000; // 5865
            16'b0001011100000011: flip_mask_bin = 48'b000000000000000000000000000000001000000000000000; // 5891
            16'b0001011101001100: flip_mask_bin = 48'b000000000000000000001101000000000000000000000000; // 5964
            16'b0001100000000000: flip_mask_bin = 48'b000110000000000000000000000000000000000000000000; // 6144
            16'b0001100111000001: flip_mask_bin = 48'b000000000000000000000000000000000000111000000000; // 6593
            16'b0001101000000000: flip_mask_bin = 48'b000110100000000000000000000000000000000000000000; // 6656
            16'b0001101011010110: flip_mask_bin = 48'b000000000000000000000000010110000000000000000000; // 6870
            16'b0001101111110111: flip_mask_bin = 48'b000000000000000000000000000000000000001010000000; // 7159
            16'b0001110000000000: flip_mask_bin = 48'b000111000000000000000000000000000000000000000000; // 7168
            16'b0001110100101110: flip_mask_bin = 48'b000000000000000000000101000000000000000000000000; // 7470
            16'b0001111000000000: flip_mask_bin = 48'b000111100000000000000000000000000000000000000000; // 7680
            16'b0001111001110110: flip_mask_bin = 48'b000000000000000010110000000000000000000000000000; // 7798
            16'b0010000000000000: flip_mask_bin = 48'b001000000000000000000000000000000000000000000000; // 8192
            16'b0010000010100011: flip_mask_bin = 48'b000000000000000000000000010010000000000000000000; // 8355
            16'b0010001110001010: flip_mask_bin = 48'b000000000000000000000000000000000000011100000000; // 9098
            16'b0010010000000000: flip_mask_bin = 48'b001001000000000000000000000000000000000000000000; // 9216
            16'b0010010011011111: flip_mask_bin = 48'b000000000000000000010100000000000000000000000000; // 9439
            16'b0010011100101011: flip_mask_bin = 48'b000000000000000000000000000000000001011000000000; // 10027
            16'b0010011111001010: flip_mask_bin = 48'b000000000000000011010000000000000000000000000000; // 10186
            16'b0010100000000000: flip_mask_bin = 48'b001010000000000000000000000000000000000000000000; // 10240
            16'b0010100000000011: flip_mask_bin = 48'b000000000000000000000000000000000011100000000000; // 10243
            16'b0010110000000000: flip_mask_bin = 48'b001011000000000000000000000000000000000000000000; // 11264
            16'b0010110101101111: flip_mask_bin = 48'b000000000000000000000001010000000000000000000000; // 11631
            16'b0010111001110100: flip_mask_bin = 48'b000000000000000000000000100000000000000000000000; // 11892
            16'b0010111001111000: flip_mask_bin = 48'b000000000000000000000000000000111000000000000000; // 11896
            16'b0010111010111101: flip_mask_bin = 48'b000000000000000000011100000000000000000000000000; // 11965
            16'b0010111100110100: flip_mask_bin = 48'b000000000000000000000000000000000000000001001000; // 12084
            16'b0010111101000101: flip_mask_bin = 48'b000000000000000000000000000001111000000000000000; // 12101
            16'b0011000000000000: flip_mask_bin = 48'b001100000000000000000000000000000000000000000000; // 12288
            16'b0011000010010111: flip_mask_bin = 48'b000000000000000000000000000000000000000000001110; // 12439
            16'b0011001101011010: flip_mask_bin = 48'b000000000000000000000101100000000000000000000000; // 13146
            16'b0011001111011110: flip_mask_bin = 48'b000000000000000001101000000000000000000000000000; // 13278
            16'b0011010000000000: flip_mask_bin = 48'b001101000000000000000000000000000000000000000000; // 13312
            16'b0011011000001111: flip_mask_bin = 48'b000000000000000000000000000000000000000000001111; // 13839
            16'b0011100000000000: flip_mask_bin = 48'b001110000000000000000000000000000000000000000000; // 14336
            16'b0011100001000110: flip_mask_bin = 48'b000000000000000000000000000001110000000000000000; // 14406
            16'b0011100001111101: flip_mask_bin = 48'b000000000000000000000000000000000000010110000000; // 14461
            16'b0011100100111011: flip_mask_bin = 48'b000000000000000000000000000000000000000000100100; // 14651
            16'b0011100101111011: flip_mask_bin = 48'b000000000000000000000000000000110000000000000000; // 14715
            16'b0011100110111100: flip_mask_bin = 48'b000000000000000001100000000000000000000000000000; // 14780
            16'b0011100110111101: flip_mask_bin = 48'b000000000000000101100000000000000000000000000000; // 14781
            16'b0011100111110010: flip_mask_bin = 48'b000000000000000000000000000000000000000000001001; // 14834
            16'b0011101001001011: flip_mask_bin = 48'b000000000000000000000000000000000000100100000000; // 14923
            16'b0011101001110101: flip_mask_bin = 48'b000000000000000000000000000100000000000000000000; // 14965
            16'b0011101101001000: flip_mask_bin = 48'b000000000000000000000000000101000000000000000000; // 15176
            16'b0011110000000000: flip_mask_bin = 48'b001111000000000000000000000000000000000000000000; // 15360
            16'b0011111011101010: flip_mask_bin = 48'b000000000000000000000000000000000001100000000000; // 16106
            16'b0011111101101010: flip_mask_bin = 48'b000000000000000000000000000000000000000000001000; // 16234
            16'b0100000000000000: flip_mask_bin = 48'b010000000000000000000000000000000000000000000000; // 16384
            16'b0100000001101011: flip_mask_bin = 48'b000000000000000000000000000000000000001110000000; // 16491
            16'b0100000111001000: flip_mask_bin = 48'b000000000000000000000000101100000000000000000000; // 16840
            16'b0100001001011101: flip_mask_bin = 48'b000000000000000000000000000000000000111100000000; // 16989
            16'b0100010110001101: flip_mask_bin = 48'b000000000000000000010110000000000000000000000000; // 17805
            16'b0100011011111100: flip_mask_bin = 48'b000000000000000000000000000000000001111000000000; // 18172
            16'b0100100000000000: flip_mask_bin = 48'b010010000000000000000000000000000000000000000000; // 18432
            16'b0100100000111110: flip_mask_bin = 48'b000000000000000000000000000000001001000000000000; // 18494
            16'b0100100100101101: flip_mask_bin = 48'b000000000000000000000000000000000000000001110000; // 18733
            16'b0100100111010100: flip_mask_bin = 48'b000000000000000000000000000000000011000000000000; // 18900
            16'b0100101111000010: flip_mask_bin = 48'b000000000000000000000000000000000000000101000000; // 19394
            16'b0100110000111101: flip_mask_bin = 48'b000000000000000000000011010000000000000000000000; // 19517
            16'b0100110011100000: flip_mask_bin = 48'b000000000000000000000000000001100000000000000000; // 19680
            16'b0100110100101010: flip_mask_bin = 48'b000000000000000000000000000000000000000011100000; // 19754
            16'b0100110111011101: flip_mask_bin = 48'b000000000000000000000000000000100000000000000000; // 19933
            16'b0100111100011111: flip_mask_bin = 48'b000000000000000000000000011110000000000000000000; // 20255
            16'b0100111100100110: flip_mask_bin = 48'b000000000000000000000010100000000000000000000000; // 20262
            16'b0100111101000000: flip_mask_bin = 48'b000000000000010110000000000000000000000000000000; // 20288
            16'b0100111101000001: flip_mask_bin = 48'b000000000000010010000000000000000000000000000000; // 20289
            16'b0100111101000010: flip_mask_bin = 48'b000000000000011110000000000000000000000000000000; // 20290
            16'b0100111101000011: flip_mask_bin = 48'b000000000000011010000000000000000000000000000000; // 20291
            16'b0100111101000100: flip_mask_bin = 48'b000000000000000110000000000000000000000000000000; // 20292
            16'b0100111101000101: flip_mask_bin = 48'b000000000000000010000000000000000000000000000000; // 20293
            16'b0100111101000110: flip_mask_bin = 48'b000000000000001110000000000000000000000000000000; // 20294
            16'b0100111101000111: flip_mask_bin = 48'b000000000000001010000000000000000000000000000000; // 20295
            16'b0100111111101111: flip_mask_bin = 48'b000000000000000000011110000000000000000000000000; // 20463
            16'b0101000000000000: flip_mask_bin = 48'b010100000000000000000000000000000000000000000000; // 20480
            16'b0101000000110101: flip_mask_bin = 48'b000000000000000000000000000000000000001111000000; // 20533
            16'b0101000011011111: flip_mask_bin = 48'b000000000000000000000000000000000000000000011010; // 20703
            16'b0101000100110011: flip_mask_bin = 48'b000000000000000000110000000000000000000000000000; // 20787
            16'b0101001000001000: flip_mask_bin = 48'b000000000000000000000111100000000000000000000000; // 21000
            16'b0101010011110100: flip_mask_bin = 48'b000000000000000000000000001001000000000000000000; // 21748
            16'b0101010111001001: flip_mask_bin = 48'b000000000000000000000000001000000000000000000000; // 21961
            16'b0101011011010010: flip_mask_bin = 48'b000000000000000000000001111000000000000000000000; // 22226
            16'b0101100000000000: flip_mask_bin = 48'b010110000000000000000000000000000000000000000000; // 22528
            16'b0101100101110011: flip_mask_bin = 48'b000000000000000000000000000000000000000000110000; // 22899
            16'b0101101011011110: flip_mask_bin = 48'b000000000000000000000000000000101000000000000000; // 23262
            16'b0101101101010001: flip_mask_bin = 48'b000000000000000000111000000000000000000000000000; // 23377
            16'b0101101110011100: flip_mask_bin = 48'b000000000000000000000000000000000000000100000000; // 23452
            16'b0101101111100011: flip_mask_bin = 48'b000000000000000000000000000001101000000000000000; // 23523
            16'b0101110101110100: flip_mask_bin = 48'b000000000000000000000000000000000000000010100000; // 23924
            16'b0101111011010111: flip_mask_bin = 48'b000000000000000000000000000000001011000000000000; // 24279
            16'b0101111100100010: flip_mask_bin = 48'b000000000000000000000000000000000000000000011100; // 24354
            16'b0101111100111101: flip_mask_bin = 48'b000000000000000000000000000000000001000000000000; // 24381
            16'b0110000000000000: flip_mask_bin = 48'b011000000000000000000000000000000000000000000000; // 24576
            16'b0110000001001000: flip_mask_bin = 48'b000000000000000000000000000000000000000000010100; // 24648
            16'b0110000101010010: flip_mask_bin = 48'b000000000000000000000010000000000000000000000000; // 24914
            16'b0110000111010111: flip_mask_bin = 48'b000000000000000000000000000000000000100000000000; // 25047
            16'b0110001001001001: flip_mask_bin = 48'b000000000000000000000011110000000000000000000000; // 25161
            16'b0110001001001111: flip_mask_bin = 48'b000000000000000000000000000000010010000000000000; // 25167
            16'b0110001010011000: flip_mask_bin = 48'b000000000000000000000000000001011000000000000000; // 25240
            16'b0110001011101101: flip_mask_bin = 48'b000000000000000001011000000000000000000000000000; // 25325
            16'b0110001110100101: flip_mask_bin = 48'b000000000000000000000000000000011000000000000000; // 25509
            16'b0110001111100001: flip_mask_bin = 48'b000000000000000000000000000000000000010010000000; // 25569
            16'b0110011000011001: flip_mask_bin = 48'b000000000000000000000000000000000000000000111000; // 26137
            16'b0110100000000000: flip_mask_bin = 48'b011010000000000000000000000000000000000000000000; // 26624
            16'b0110100010001111: flip_mask_bin = 48'b000000000000000001010000000000000000000000000000; // 26767
            16'b0110101100110000: flip_mask_bin = 48'b000000000000000000001010000000000000000000000000; // 27440
            16'b0110111010000001: flip_mask_bin = 48'b000000000000000000000000001101000000000000000000; // 28289
            16'b0110111110110101: flip_mask_bin = 48'b000000000000000000000000000000000000000000010010; // 28597
            16'b0110111110111100: flip_mask_bin = 48'b000000000000000000000000001100000000000000000000; // 28604
            16'b0111000000000000: flip_mask_bin = 48'b011100000000000000000000000000000000000000000000; // 28672
            16'b0111010010100110: flip_mask_bin = 48'b000000000000000000000000000000010000000000000000; // 29862
            16'b0111010101001100: flip_mask_bin = 48'b000000000000000000000000000000011010000000000000; // 30028
            16'b0111010101101010: flip_mask_bin = 48'b000000000000000000000000011010000000000000000000; // 30058
            16'b0111010110011011: flip_mask_bin = 48'b000000000000000000000000000001010000000000000000; // 30107
            16'b0111010111101100: flip_mask_bin = 48'b000000000000000000100100000000000000000000000000; // 30188
            16'b0111011000011110: flip_mask_bin = 48'b000000000000000000001111000000000000000000000000; // 30238
            16'b0111011001000111: flip_mask_bin = 48'b000000000000000000000000000000000000000001111000; // 30279
            16'b0111011010010101: flip_mask_bin = 48'b000000000000000000000000000101100000000000000000; // 30357
            16'b0111011011111000: flip_mask_bin = 48'b000000000000000111100000000000000000000000000000; // 30456
            16'b0111011011111001: flip_mask_bin = 48'b000000000000000011100000000000000000000000000000; // 30457
            16'b0111011100111110: flip_mask_bin = 48'b000000000000000000000000000000000010100000000000; // 30526
            16'b0111011110101000: flip_mask_bin = 48'b000000000000000000000000000100100000000000000000; // 30632
            16'b0111100000000000: flip_mask_bin = 48'b011110000000000000000000000000000000000000000000; // 30720
            16'b0111100000010110: flip_mask_bin = 48'b000000000000000000000000000000000000011000000000; // 30742
            16'b0111100010100110: flip_mask_bin = 48'b000000000000000000000001011000000000000000000000; // 30886
            16'b0111101110111101: flip_mask_bin = 48'b000000000000000000000000101000000000000000000000; // 31677
            16'b0111110001111100: flip_mask_bin = 48'b000000000000000000000111000000000000000000000000; // 31868
            16'b0111111110001110: flip_mask_bin = 48'b000000000000000000101100000000000000000000000000; // 32654
            16'b1000000000000000: flip_mask_bin = 48'b100000000000000000000000000000000000000000000000; // 32768
            16'b1000001000111001: flip_mask_bin = 48'b000000000000000010010000000000000000000000000000; // 33337
            16'b1000001010010011: flip_mask_bin = 48'b000000000000000000001110000000000000000000000000; // 33427
            16'b1000010010110001: flip_mask_bin = 48'b000000000000000000000000000000000011010000000000; // 33969
            16'b1000010110110111: flip_mask_bin = 48'b000000000000000000000000000000000000000001011000; // 34231
            16'b1000100011110001: flip_mask_bin = 48'b000000000000000000000110000000000000000000000000; // 35057
            16'b1000101110011001: flip_mask_bin = 48'b000000000000000000000000000000000001101000000000; // 35737
            16'b1000110000101011: flip_mask_bin = 48'b000000000000000000000000011000000000000000000000; // 35883
            16'b1000110011011010: flip_mask_bin = 48'b000000000000000000000000000011010000000000000000; // 36058
            16'b1000110100001110: flip_mask_bin = 48'b000000000000000000000000000000000000011110000000; // 36110
            16'b1000110111100111: flip_mask_bin = 48'b000000000000000000000000000010010000000000000000; // 36327
            16'b1000111001110010: flip_mask_bin = 48'b000000000000000000000000000000001100000000000000; // 36466
            16'b1000111011101001: flip_mask_bin = 48'b000000000000000000000000000110100000000000000000; // 36585
            16'b1000111100110000: flip_mask_bin = 48'b000000000000000000000001101000000000000000000000; // 36656
            16'b1000111100111000: flip_mask_bin = 48'b000000000000000000000000000000000000101100000000; // 36664
            16'b1000111110011000: flip_mask_bin = 48'b000000000000000000000000000000000110000000000000; // 36760
            16'b1000111111010100: flip_mask_bin = 48'b000000000000000000000000000111100000000000000000; // 36820
            16'b1001000000000000: flip_mask_bin = 48'b100100000000000000000000000000000000000000000000; // 36864
            16'b1001001001011000: flip_mask_bin = 48'b000000000000000000000000000000000001010000000000; // 37464
            16'b1001001110111000: flip_mask_bin = 48'b000000000000000000000000000000000000000000110100; // 37816
            16'b1001010111011111: flip_mask_bin = 48'b000000000000000000000011000000000000000000000000; // 38367
            16'b1001010111101001: flip_mask_bin = 48'b000000000000000000000000000000000000000000011000; // 38377
            16'b1001011000101101: flip_mask_bin = 48'b000000000000000000101000000000000000000000000000; // 38445
            16'b1001011011000100: flip_mask_bin = 48'b000000000000000000000010110000000000000000000000; // 38596
            16'b1001011011111001: flip_mask_bin = 48'b000000000000000000000000000000000000010100000000; // 38649
            16'b1001011011111101: flip_mask_bin = 48'b000000000000000000000000001110000000000000000000; // 38653
            16'b1001011111000000: flip_mask_bin = 48'b000000000000000000000000001111000000000000000000; // 38848
            16'b1001100000101010: flip_mask_bin = 48'b000000000000000000000000111100000000000000000000; // 38954
            16'b1001100010011011: flip_mask_bin = 48'b000000000000000000000000000000001110000000000000; // 39067
            16'b1001100101110001: flip_mask_bin = 48'b000000000000000000000000000000000100000000000000; // 39281
            16'b1001101000010100: flip_mask_bin = 48'b000000000000000000000000000000000000000000011110; // 39444
            16'b1001110001001110: flip_mask_bin = 48'b000000000000000100100000000000000000000000000000; // 40014
            16'b1001110001001111: flip_mask_bin = 48'b000000000000000000100000000000000000000000000000; // 40015
            16'b1001111110111101: flip_mask_bin = 48'b000000000000000000001011000000000000000000000000; // 40893
            16'b1010000000000000: flip_mask_bin = 48'b101000000000000000000000000000000000000000000000; // 40960
            16'b1010000000001010: flip_mask_bin = 48'b000000000000000000000000000000110100000000000000; // 40970
            16'b1010000101000100: flip_mask_bin = 48'b000000000000000000000001001000000000000000000000; // 41284
            16'b1010001001011111: flip_mask_bin = 48'b000000000000000000000000111000000000000000000000; // 41567
            16'b1010010100101101: flip_mask_bin = 48'b000000000000000000000000000000000000001001000000; // 42285
            16'b1010010101111110: flip_mask_bin = 48'b000000000000000000000000000000000000000000010110; // 42366
            16'b1010010111110000: flip_mask_bin = 48'b000000000000001101000000000000000000000000000000; // 42480
            16'b1010010111110001: flip_mask_bin = 48'b000000000000001001000000000000000000000000000000; // 42481
            16'b1010010111110010: flip_mask_bin = 48'b000000000000000101000000000000000000000000000000; // 42482
            16'b1010010111110011: flip_mask_bin = 48'b000000000000000001000000000000000000000000000000; // 42483
            16'b1010011001001100: flip_mask_bin = 48'b000000000000000000011010000000000000000000000000; // 42572
            16'b1010011010000101: flip_mask_bin = 48'b000000000000000000000110100000000000000000000000; // 42629
            16'b1010011110011011: flip_mask_bin = 48'b000000000000000000000000000000000101100000000000; // 42907
            16'b1010100001101100: flip_mask_bin = 48'b000000000000000000000000000000000000000100100000; // 43116
            16'b1010101010000011: flip_mask_bin = 48'b000000000000000000000000000000000000000000010000; // 43651
            16'b1010110000101110: flip_mask_bin = 48'b000000000000000000010010000000000000000000000000; // 44078
            16'b1010110010001000: flip_mask_bin = 48'b000000000000000000000000001010000000000000000000; // 44168
            16'b1010110010110010: flip_mask_bin = 48'b000000000000000000000000000000000000110000000000; // 44210
            16'b1010110011010010: flip_mask_bin = 48'b000000000000000000000000000000000000000000111100; // 44242
            16'b1010110110110101: flip_mask_bin = 48'b000000000000000000000000001011000000000000000000; // 44469
            16'b1010111010000100: flip_mask_bin = 48'b000000000000000000000000000000000000000010000000; // 44676
            16'b1010111110010001: flip_mask_bin = 48'b000000000000000001001000000000000000000000000000; // 44945
            16'b1011000000000000: flip_mask_bin = 48'b101100000000000000000000000000000000000000000000; // 45056
            16'b1011000101110010: flip_mask_bin = 48'b000000000000000000000000000000000111100000000000; // 45426
            16'b1011001011110010: flip_mask_bin = 48'b000000000000000000111100000000000000000000000000; // 45810
            16'b1011010010011100: flip_mask_bin = 48'b000000000000000000000000000010100000000000000000; // 46236
            16'b1011010101110011: flip_mask_bin = 48'b000000000000000000000000000000000000001000000000; // 46451
            16'b1011010110100001: flip_mask_bin = 48'b000000000000000000000000000011100000000000000000; // 46497
            16'b1011011001011110: flip_mask_bin = 48'b000000000000000000000000011100000000000000000000; // 46686
            16'b1011011100001001: flip_mask_bin = 48'b000000000000000000000000000000111100000000000000; // 46857
            16'b1011100000110010: flip_mask_bin = 48'b000000000000000000000000000000000000000101100000; // 47154
            16'b1011100010010000: flip_mask_bin = 48'b000000000000000000110100000000000000000000000000; // 47248
            16'b1011100010110000: flip_mask_bin = 48'b000000000000000000000010010000000000000000000000; // 47280
            16'b1011101001011011: flip_mask_bin = 48'b000000000000000000000000000000000010110000000000; // 47707
            16'b1011101011011101: flip_mask_bin = 48'b000000000000000000000000000000000000000001010000; // 47837
            16'b1011101110000101: flip_mask_bin = 48'b000000000000000011110000000000000000000000000000; // 48005
            16'b1011101110101011: flip_mask_bin = 48'b000000000000000000000011100000000000000000000000; // 48043
            16'b1011111011011010: flip_mask_bin = 48'b000000000000000000000000000000000000000011000000; // 48858
            16'b1100000000000000: flip_mask_bin = 48'b110000000000000000000000000000000000000000000000; // 49152
            16'b1100000000111010: flip_mask_bin = 48'b000000000000000000000000000010110000000000000000; // 49210
            16'b1100000100000111: flip_mask_bin = 48'b000000000000000000000000000011110000000000000000; // 49415
            16'b1100001000001001: flip_mask_bin = 48'b000000000000000000000000000111000000000000000000; // 49673
            16'b1100001100110100: flip_mask_bin = 48'b000000000000000000000000000110000000000000000000; // 49972
            16'b1100001110101110: flip_mask_bin = 48'b000000000000000000000000000000000000000000000011; // 50094
            16'b1100001110101111: flip_mask_bin = 48'b000000000000000000000000000000101100000000000000; // 50095
            16'b1100010100110110: flip_mask_bin = 48'b000000000000000000000000000000000000000000000010; // 50486
            16'b1100011001001100: flip_mask_bin = 48'b000000000000000000000000000000000101000000000000; // 50764
            16'b1100011100011110: flip_mask_bin = 48'b000000000000000000011000000000000000000000000000; // 50974
            16'b1100011110100110: flip_mask_bin = 48'b000000000000000000000000000000001111000000000000; // 51110
            16'b1100011111010111: flip_mask_bin = 48'b000000000000000000000100100000000000000000000000; // 51159
            16'b1100101011001011: flip_mask_bin = 48'b000000000000000000000000000000000000000000000100; // 51915
            16'b1100110001010011: flip_mask_bin = 48'b000000000000000000000000000000000000000000000101; // 52307
            16'b1100110010011010: flip_mask_bin = 48'b000000000000000000000000000000000000000000101000; // 52378
            16'b1100110101100101: flip_mask_bin = 48'b000000000000000000000000000000000000010000000000; // 52581
            16'b1100110101111100: flip_mask_bin = 48'b000000000000000000010000000000000000000000000000; // 52604
            16'b1100110111100011: flip_mask_bin = 48'b000000000000000000000000110100000000000000000000; // 52707
            16'b1101000000000000: flip_mask_bin = 48'b110100000000000000000000000000000000000000000000; // 53248
            16'b1101000010100101: flip_mask_bin = 48'b000000000000000000000000000000000111000000000000; // 53413
            16'b1101000101001111: flip_mask_bin = 48'b000000000000000000000000000000001101000000000000; // 53583
            16'b1101001100001010: flip_mask_bin = 48'b000000000000000010100000000000000000000000000000; // 54026
            16'b1101001100001011: flip_mask_bin = 48'b000000000000000110100000000000000000000000000000; // 54027
            16'b1101010010100100: flip_mask_bin = 48'b000000000000000000000000000000000000101000000000; // 54436
            16'b1101010010101100: flip_mask_bin = 48'b000000000000000000000000000000100100000000000000; // 54444
            16'b1101011010010010: flip_mask_bin = 48'b000000000000000000000000000000000000011010000000; // 54930
            16'b1101100111100010: flip_mask_bin = 48'b000000000000000000000000010000000000000000000000; // 55778
            16'b1101101011111001: flip_mask_bin = 48'b000000000000000000000001100000000000000000000000; // 56057
            16'b1101101110001100: flip_mask_bin = 48'b000000000000000000000000000000000010010000000000; // 56204
            16'b1101110011000100: flip_mask_bin = 48'b000000000000000000000000000000000000000001101000; // 56516
            16'b1110000000000000: flip_mask_bin = 48'b111000000000000000000000000000000000000000000000; // 57344
            16'b1110001110010111: flip_mask_bin = 48'b000000000000000000000000010100000000000000000000; // 58263
            16'b1110001110101110: flip_mask_bin = 48'b000000000000000000000000000000000000000001100000; // 58286
            16'b1110001111000001: flip_mask_bin = 48'b000000000000000000001100000000000000000000000000; // 58305
            16'b1110010101000110: flip_mask_bin = 48'b000000000000000000000000000000000000000111000000; // 58694
            16'b1110010101100110: flip_mask_bin = 48'b000000000000000000000000000000000011110000000000; // 58726
            16'b1110011110101001: flip_mask_bin = 48'b000000000000000000000000000000000000000011110000; // 59305
            16'b1110100110100011: flip_mask_bin = 48'b000000000000000000000100000000000000000000000000; // 59811
            16'b1110101001001110: flip_mask_bin = 48'b000000000000000000000000000000000001001000000000; // 59982
            16'b1110101010110100: flip_mask_bin = 48'b000000000000001011000000000000000000000000000000; // 60084
            16'b1110101010110101: flip_mask_bin = 48'b000000000000001111000000000000000000000000000000; // 60085
            16'b1110101010110110: flip_mask_bin = 48'b000000000000000011000000000000000000000000000000; // 60086
            16'b1110101010110111: flip_mask_bin = 48'b000000000000000111000000000000000000000000000000; // 60087
            16'b1110110000111101: flip_mask_bin = 48'b000000000000000000000000000000011110000000000000; // 60477
            16'b1110110111010111: flip_mask_bin = 48'b000000000000000000000000000000010100000000000000; // 60887
            16'b1110111001001111: flip_mask_bin = 48'b000000000000000000000000000000000110100000000000; // 61007
            16'b1110111011101111: flip_mask_bin = 48'b000000000000000000000000000000000000001100000000; // 61167
            16'b1111000000000000: flip_mask_bin = 48'b111100000000000000000000000000000000000000000000; // 61440
            16'b1111001100111001: flip_mask_bin = 48'b000000000000000000000000000000000000000000001101; // 62265
            16'b1111001110001111: flip_mask_bin = 48'b000000000000000000000000000000000001110000000000; // 62351
            16'b1111001111110000: flip_mask_bin = 48'b000000000000000000000000000000000000000000100000; // 62448
            16'b1111010010001101: flip_mask_bin = 48'b000000000000000000000001000000000000000000000000; // 62605
            16'b1111010011000000: flip_mask_bin = 48'b000000000000000001110000000000000000000000000000; // 62656
            16'b1111010100011000: flip_mask_bin = 48'b000000000000000000000000000000000000000110000000; // 62744
            16'b1111010110100001: flip_mask_bin = 48'b000000000000000000000000000000000000000000001100; // 62881
            16'b1111011100101110: flip_mask_bin = 48'b000000000000000000000000000000000000110100000000; // 63278
            16'b1111011110010110: flip_mask_bin = 48'b000000000000000000000000110000000000000000000000; // 63382
            16'b1111011111110111: flip_mask_bin = 48'b000000000000000000000000000000000000000010110000; // 63479
            16'b1111100001111100: flip_mask_bin = 48'b000000000000000000000000000011000000000000000000; // 63612
            16'b1111100010100110: flip_mask_bin = 48'b000000000000000000000000000000000100100000000000; // 63654
            16'b1111100101000001: flip_mask_bin = 48'b000000000000000000000000000010000000000000000000; // 63809
            16'b1111101001011100: flip_mask_bin = 48'b000000000000000001111000000000000000000000000000; // 64092
            16'b1111101011010100: flip_mask_bin = 48'b000000000000000000000000000000011100000000000000; // 64212
            16'b1111101100111110: flip_mask_bin = 48'b000000000000000000000000000000010110000000000000; // 64318
            16'b1111110011000100: flip_mask_bin = 48'b000000000000000000000000000000000000000000001011; // 64708
            16'b1111111010100010: flip_mask_bin = 48'b000000000000000001111000000000000000000000000000; // 65186
            16'b1111111010110001: flip_mask_bin = 48'b000000000000000000000000000000000000001101000000; // 65201
            16'b1111111011101111: flip_mask_bin = 48'b000000000000000000001001000000000000000000000000; // 65263
            default: flip_mask_bin = 48'b0;
        endcase
    end
endmodule
